--freq_demod test
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity freq_demod_test is
	--
end freq_demod_test;

architecture sim of freq_demod_test is
	component freq_demod is
		port(
			clk_i		: in std_logic;									-- demod clock
			i_i, q_i	: in signed(15 downto 0);						-- I/Q inputs
			demod_o		: out signed(15 downto 0) := (others => '0')	-- freq demod out
		);
	end component;

	signal clk_i : std_logic := '0';
	signal i_i, q_i, demod_o : signed(15 downto 0) := (others => '0');

	type vals is array(0 to 20000-1) of signed(15 downto 0);
	constant i_vals : vals := (
		x"FB53", x"F825", x"F463", x"F0C4", x"EDC8", x"EC13", x"EBF3", x"EDB9",
		x"F195", x"F77E", x"FEE8", x"069F", x"0D49", x"11DF", x"13B2", x"1284",
		x"0EBB", x"0928", x"0297", x"FB9A", x"F4ED", x"EF9A", x"ECA0", x"ED42",
		x"F18F", x"F89F", x"009D", x"07F2", x"0DA5", x"113D", x"127D", x"11BF",
		x"0F74", x"0C7C", x"095D", x"068D", x"0488", x"03D3", x"04F7", x"07E9",
		x"0BF9", x"1016", x"12FA", x"1348", x"1062", x"0A36", x"01E3", x"F8EB",
		x"F184", x"ED3E", x"ECD7", x"EF93", x"F3F3", x"F856", x"FB2B", x"FB5A",
		x"F8AE", x"F452", x"EFF8", x"ED5A", x"EDB5", x"F136", x"F714", x"FE0C",
		x"0490", x"0993", x"0CD7", x"0ECE", x"0FB4", x"0FFC", x"0FF6", x"0FDE",
		x"0FDC", x"0FC6", x"0F50", x"0E82", x"0D1D", x"0AB4", x"06CC", x"014E",
		x"FABD", x"F43B", x"EF29", x"EC7E", x"ECC5", x"EFAA", x"F412", x"F8BE",
		x"FC89", x"FF02", x"FFCF", x"FF19", x"FD00", x"F9BD", x"F5D0", x"F1F2",
		x"EEB5", x"ECF8", x"ED5B", x"F078", x"F63E", x"FDD7", x"058D", x"0BD8",
		x"0FDF", x"119A", x"116B", x"0FAD", x"0CDB", x"0934", x"054C", x"023A",
		x"0122", x"02BD", x"06B2", x"0BE5", x"108A", x"12C3", x"11AF", x"0DCB",
		x"089D", x"03D9", x"00A1", x"FF4E", x"FFF4", x"0269", x"0612", x"0A17",
		x"0E13", x"115A", x"1397", x"143C", x"12B0", x"0EA5", x"0876", x"0109",
		x"F99D", x"F352", x"EEE4", x"EC41", x"EB19", x"EACA", x"EB05", x"EB5A",
		x"EBD1", x"EC61", x"ED0E", x"EE15", x"EFA6", x"F1ED", x"F46E", x"F6F6",
		x"F95A", x"FBCE", x"FE16", x"0060", x"0272", x"0467", x"065F", x"0898",
		x"0B25", x"0DD2", x"106F", x"12B5", x"143E", x"1465", x"1246", x"0D97",
		x"06B1", x"FE93", x"F6B6", x"F071", x"ECCB", x"EC08", x"EDFF", x"F236",
		x"F7E8", x"FEA5", x"05D1", x"0C8E", x"1146", x"12BB", x"102C", x"0A4E",
		x"02BC", x"FB62", x"F593", x"F228", x"F16C", x"F354", x"F788", x"FD66",
		x"044D", x"0B0C", x"1065", x"1298", x"10B7", x"0AD6", x"0241", x"F920",
		x"F19E", x"ECFC", x"EB5C", x"EB5A", x"EB86", x"EB8E", x"EB9C", x"ECF4",
		x"F0A5", x"F6EA", x"FEFB", x"06E8", x"0CE7", x"0F67", x"0E24", x"096A",
		x"0260", x"FA4B", x"F2F2", x"EE0D", x"EC59", x"EDA0", x"F092", x"F39F",
		x"F5D0", x"F71A", x"F7DF", x"F919", x"FB7F", x"FFAC", x"052F", x"0B42",
		x"1053", x"1318", x"12F8", x"0FD6", x"0A8B", x"0480", x"FED5", x"FA11",
		x"F679", x"F3B8", x"F191", x"EFE3", x"EE7E", x"ED64", x"EC86", x"EBF8",
		x"EB77", x"EAFC", x"EA8B", x"EA53", x"EAB2", x"EBF7", x"EE61", x"F2A2",
		x"F8F9", x"0109", x"0938", x"0F99", x"134A", x"1494", x"148C", x"144F",
		x"145B", x"1474", x"1388", x"104D", x"09FE", x"015B", x"F879", x"F171",
		x"ED4B", x"EC21", x"EDB3", x"F16C", x"F6DF", x"FD73", x"04A7", x"0BA4",
		x"1101", x"130F", x"10E6", x"0B4F", x"03C4", x"FC59", x"F63D", x"F279",
		x"F1DD", x"F4C8", x"FAC8", x"028B", x"0A2F", x"0FEF", x"130C", x"13A3",
		x"1271", x"111F", x"10BE", x"117C", x"12DB", x"1433", x"14CA", x"14DB",
		x"14B7", x"146C", x"13E5", x"126D", x"0EF3", x"0915", x"0139", x"F8F7",
		x"F203", x"EDBD", x"ECAA", x"EED1", x"F3C5", x"FA88", x"01EB", x"08BE",
		x"0E29", x"11DD", x"13EE", x"14CB", x"14F3", x"14B7", x"142D", x"136D",
		x"127B", x"114D", x"0FAA", x"0D67", x"0A7C", x"0761", x"0456", x"01BF",
		x"FFD9", x"FEA5", x"FE5E", x"FEC2", x"FFD6", x"0142", x"02DD", x"04DC",
		x"0796", x"0B59", x"0F87", x"12B2", x"1378", x"10E0", x"0B56", x"03F7",
		x"FC37", x"F5EB", x"F273", x"F2EF", x"F786", x"FEFF", x"0740", x"0DFA",
		x"1212", x"137B", x"1393", x"1379", x"13B4", x"13CA", x"1279", x"0EE3",
		x"0864", x"0044", x"F88C", x"F2EB", x"F016", x"EF7E", x"F027", x"F1AD",
		x"F42A", x"F7E9", x"FCD4", x"029F", x"08A9", x"0E15", x"11D1", x"12F7",
		x"111D", x"0CAB", x"06F0", x"018B", x"FDE6", x"FC96", x"FD6C", x"FFC7",
		x"0312", x"06C0", x"0A69", x"0D38", x"0EFA", x"0F2B", x"0E6E", x"0CB3",
		x"0A7E", x"07C4", x"0492", x"010F", x"FD5C", x"F9B1", x"F633", x"F2FD",
		x"F02C", x"EDF6", x"EC85", x"EBE0", x"EBF2", x"ED0D", x"EF9F", x"F42D",
		x"FACA", x"027D", x"0A28", x"103D", x"13AF", x"142D", x"12C3", x"108B",
		x"0E96", x"0D3E", x"0C58", x"0B4B", x"09C6", x"0765", x"0416", x"0041",
		x"FC26", x"F80E", x"F4A1", x"F209", x"F116", x"F1B0", x"F3F5", x"F824",
		x"FE0D", x"04F0", x"0BB3", x"10EB", x"13A5", x"1388", x"10D7", x"0C84",
		x"0753", x"0285", x"FE87", x"FBCC", x"FA9F", x"FAE3", x"FC9E", x"FFB6",
		x"040F", x"092B", x"0E5E", x"1259", x"13E3", x"120F", x"0CB7", x"0492",
		x"FB7C", x"F368", x"EE12", x"EBE5", x"ECDC", x"EFD2", x"F38D", x"F685",
		x"F7BA", x"F6FC", x"F4D0", x"F210", x"EF55", x"ED33", x"EBF3", x"EB86",
		x"EC98", x"EF87", x"F485", x"FB82", x"038A", x"0B48", x"115A", x"148C",
		x"14E9", x"137F", x"11AA", x"1061", x"0FA5", x"0EE9", x"0D56", x"0A90",
		x"0618", x"FFF2", x"F8DE", x"F27D", x"EDF7", x"EC90", x"EDFE", x"F12C",
		x"F4B1", x"F705", x"F7A9", x"F69B", x"F458", x"F1C5", x"EF5A", x"ED9A",
		x"EC6D", x"EBCC", x"EB87", x"EBAF", x"EC7A", x"EDAF", x"EF83", x"F20E",
		x"F5B4", x"FAA3", x"0063", x"0681", x"0C51", x"10E7", x"138D", x"1373",
		x"1044", x"0A44", x"0272", x"FA5B", x"F338", x"EE2B", x"EBC6", x"EC16",
		x"EEA5", x"F2C3", x"F798", x"FC6B", x"008D", x"03C5", x"0610", x"07B6",
		x"091A", x"0AA6", x"0CAD", x"0EEF", x"1133", x"1301", x"1451", x"1500",
		x"1557", x"1575", x"155D", x"1490", x"123F", x"0D8E", x"06B2", x"FE7D",
		x"F66A", x"F007", x"EC16", x"EB43", x"ED9E", x"F2F2", x"FA80", x"02BD",
		x"0A6C", x"1092", x"1490", x"1633", x"1583", x"127F", x"0D48", x"0664",
		x"FE41", x"F624", x"EF64", x"EB63", x"EAB1", x"ED6C", x"F2F4", x"FA6C",
		x"02B8", x"0A85", x"1096", x"143C", x"159B", x"15A2", x"1531", x"14CB",
		x"140C", x"129D", x"10DF", x"0F37", x"0E49", x"0E4C", x"0F5B", x"10E9",
		x"1293", x"13D8", x"14AE", x"1528", x"155C", x"156E", x"1547", x"14F4",
		x"1466", x"13A7", x"129B", x"111A", x"0F03", x"0C86", x"09E1", x"0761",
		x"052B", x"0324", x"00F8", x"FE78", x"FBD5", x"F909", x"F60E", x"F323",
		x"F06B", x"EE2A", x"ECA1", x"EBC4", x"EB4E", x"EB25", x"EB4E", x"EBB7",
		x"EC9B", x"EDE2", x"EF79", x"F15D", x"F30F", x"F47C", x"F561", x"F5B6",
		x"F555", x"F430", x"F281", x"F058", x"EE35", x"EC83", x"EBC3", x"EC6F",
		x"EEE0", x"F350", x"F967", x"00B0", x"0826", x"0EA8", x"12D0", x"13D4",
		x"1161", x"0BFA", x"04A3", x"FCCC", x"F5B1", x"F048", x"ECCA", x"EB02",
		x"EA99", x"EB2D", x"EC6F", x"EDE7", x"EF46", x"F0A1", x"F205", x"F3A3",
		x"F538", x"F6D8", x"F8AD", x"FA99", x"FCA5", x"FF1B", x"0283", x"0705",
		x"0C3F", x"10B9", x"12D7", x"11AA", x"0D45", x"06C1", x"002A", x"FB65",
		x"FA4F", x"FD65", x"03AA", x"0ACF", x"103C", x"1256", x"118A", x"0F4B",
		x"0D93", x"0DBD", x"0FA0", x"11AB", x"1178", x"0D71", x"0680", x"FEEE",
		x"FA0C", x"F9CC", x"FE2E", x"056E", x"0CD6", x"11C0", x"1311", x"11C7",
		x"0FAE", x"0E93", x"0F5B", x"1150", x"12C7", x"11AD", x"0D3A", x"0647",
		x"FEF2", x"F957", x"F673", x"F66E", x"F8A5", x"FC75", x"00BB", x"04BE",
		x"07E6", x"09E1", x"0A6D", x"09AD", x"07B8", x"050B", x"01DC", x"FE80",
		x"FB06", x"F7C5", x"F50E", x"F2E8", x"F128", x"EF95", x"EE1D", x"ECB2",
		x"EB89", x"EAA1", x"EA26", x"EA69", x"EB41", x"EC4D", x"ED61", x"EE79",
		x"EFD8", x"F1B8", x"F3F8", x"F67F", x"F97D", x"FCDF", x"008D", x"0418",
		x"0702", x"08F5", x"09B9", x"0950", x"07EC", x"0575", x"022C", x"FE69",
		x"FADB", x"F839", x"F71E", x"F7F7", x"FAD9", x"FFC2", x"05F9", x"0C44",
		x"1107", x"132E", x"11FA", x"0D61", x"0677", x"FE94", x"F737", x"F164",
		x"ED7E", x"EBF9", x"ED07", x"F0CA", x"F6BC", x"FE3C", x"0643", x"0D52",
		x"1219", x"13F6", x"1316", x"1033", x"0C43", x"07E2", x"0407", x"00D3",
		x"FE89", x"FCAF", x"FAEE", x"F902", x"F6B5", x"F421", x"F15A", x"EEAF",
		x"ECA0", x"EB70", x"EAFC", x"EAB1", x"EA72", x"EAC1", x"ECB8", x"F133",
		x"F817", x"002D", x"07EB", x"0E60", x"12CC", x"14F8", x"14FF", x"1303",
		x"0F18", x"0907", x"013C", x"F895", x"F155", x"ED66", x"EDB6", x"F231",
		x"F9B0", x"0269", x"0A4D", x"103C", x"13E8", x"15C1", x"15F4", x"148F",
		x"113E", x"0BBC", x"043F", x"FBBF", x"F3D9", x"EE0A", x"EAE9", x"E9EE",
		x"EA5A", x"EB8A", x"ED4F", x"EFAA", x"F283", x"F526", x"F6DD", x"F6FB",
		x"F557", x"F2AD", x"EFCC", x"ED67", x"EBDD", x"EB07", x"EADF", x"EB85",
		x"EDA3", x"F1B0", x"F7E2", x"FF8B", x"0765", x"0E0D", x"128F", x"1496",
		x"1484", x"1329", x"1169", x"0FB4", x"0E41", x"0CF1", x"0BA6", x"0A32",
		x"080B", x"0506", x"0162", x"FDBA", x"FA4B", x"F758", x"F4F2", x"F386",
		x"F372", x"F4B1", x"F6EC", x"FA39", x"FDF7", x"01B9", x"04CE", x"06A9",
		x"0703", x"05EA", x"03AB", x"005F", x"FCB7", x"F919", x"F657", x"F4F7",
		x"F521", x"F72F", x"FB03", x"0061", x"06DB", x"0D26", x"11D9", x"137A",
		x"113D", x"0B90", x"038A", x"FB07", x"F3A1", x"EE7D", x"EC0E", x"EC01",
		x"EDB4", x"EFC0", x"F13E", x"F1B7", x"F106", x"EF66", x"ED87", x"EBEC",
		x"EB1A", x"EB2C", x"EBC3", x"ECBB", x"EE0D", x"EF5B", x"F096", x"F1E2",
		x"F392", x"F5B3", x"F878", x"FBFE", x"0019", x"043B", x"082D", x"0B24",
		x"0CF7", x"0D5E", x"0BED", x"0843", x"0266", x"FB29", x"F423", x"EF20",
		x"ECFB", x"ED6F", x"EF0B", x"F078", x"F0A8", x"EFB4", x"EDF0", x"EC37",
		x"EB46", x"EAFD", x"EAF0", x"EB16", x"EC41", x"EF91", x"F592", x"FD7A",
		x"05A6", x"0CAD", x"1199", x"13C6", x"135B", x"103A", x"0AD7", x"03A8",
		x"FB92", x"F3FA", x"EE57", x"EBA6", x"EBEC", x"EDF8", x"F098", x"F2DE",
		x"F487", x"F5A8", x"F69E", x"F75C", x"F796", x"F72F", x"F600", x"F462",
		x"F26D", x"F076", x"EE9C", x"ED1B", x"EBFB", x"EB36", x"EADB", x"EB03",
		x"EB42", x"EBE5", x"ECB2", x"EDF2", x"EFD6", x"F27B", x"F5C0", x"F952",
		x"FD1E", x"00B5", x"03B7", x"0559", x"052B", x"02C0", x"FE11", x"F7CA",
		x"F19A", x"ED6A", x"EC99", x"EEF8", x"F2EA", x"F6A9", x"F8B2", x"F881",
		x"F66A", x"F336", x"F018", x"EDB5", x"EC51", x"EBE0", x"ECE7", x"EF7C",
		x"F3EF", x"FA47", x"01FE", x"09FA", x"105B", x"1383", x"129F", x"0E60",
		x"07D6", x"0046", x"F8EE", x"F2AD", x"EE2F", x"EBDA", x"EBB7", x"ED23",
		x"EF71", x"F215", x"F483", x"F68D", x"F806", x"F8D6", x"F90E", x"F8B0",
		x"F7D8", x"F63E", x"F458", x"F211", x"EFE4", x"EDF3", x"EC5C", x"EB41",
		x"EAD1", x"EAC7", x"EAE8", x"EB15", x"EB52", x"EC1B", x"EDC7", x"F0F6",
		x"F638", x"FDB5", x"0637", x"0DBD", x"1276", x"1415", x"13AB", x"12E2",
		x"12DE", x"135D", x"1325", x"10F9", x"0BF0", x"0495", x"FC70", x"F59E",
		x"F198", x"F0B1", x"F21D", x"F50D", x"F8D1", x"FD02", x"00AF", x"02D7",
		x"027F", x"FFAD", x"FB0C", x"F580", x"F071", x"ED75", x"ED97", x"F10D",
		x"F781", x"FF88", x"07D8", x"0EA1", x"12A0", x"1374", x"1170", x"0DDB",
		x"09FF", x"0740", x"0630", x"071E", x"0984", x"0CA0", x"0FBC", x"121B",
		x"13AB", x"145A", x"145D", x"1385", x"11D7", x"0F86", x"0CBF", x"0A12",
		x"07CE", x"0640", x"05A5", x"05D1", x"06B0", x"081C", x"09FD", x"0C74",
		x"0F34", x"1213", x"13F9", x"141F", x"118E", x"0C4C", x"051B", x"FD33",
		x"F601", x"F084", x"ED5F", x"EC70", x"ECEC", x"EE3D", x"F04B", x"F309",
		x"F628", x"F94D", x"FB5D", x"FBDC", x"FAAB", x"F82F", x"F52E", x"F259",
		x"F006", x"EE5F", x"ED66", x"ECD4", x"ECC5", x"ED22", x"EDF3", x"EEF7",
		x"F0AF", x"F37F", x"F7B8", x"FD49", x"03E7", x"0AA8", x"103C", x"1373",
		x"13CB", x"1175", x"0D58", x"08FC", x"05A1", x"03DD", x"03F2", x"0599",
		x"0855", x"0BD7", x"0F5B", x"1250", x"142B", x"1513", x"1532", x"14F0",
		x"1490", x"13FE", x"1374", x"12FC", x"12A2", x"1276", x"1288", x"12C5",
		x"1357", x"143C", x"14F9", x"151D", x"13E4", x"1073", x"0ACD", x"0362",
		x"FB62", x"F431", x"EECA", x"EBCA", x"EAD0", x"EB46", x"EC1E", x"ECA4",
		x"ECA0", x"EC1E", x"EBA0", x"EB96", x"ECC3", x"EF9E", x"F4B2", x"FBBB",
		x"03AE", x"0B10", x"107C", x"1365", x"1438", x"139B", x"1294", x"11B3",
		x"1174", x"1230", x"138E", x"14A6", x"147B", x"128D", x"0FC0", x"0DE0",
		x"0E5A", x"10B3", x"12DB", x"12B6", x"0FC1", x"0B22", x"06A6", x"035E",
		x"01A5", x"017C", x"0336", x"0680", x"0AD8", x"0F15", x"129E", x"1476",
		x"1439", x"11AD", x"0CCD", x"061E", x"FEBE", x"F781", x"F1B9", x"EDE1",
		x"EBDC", x"EB04", x"EAC2", x"EAF1", x"EB3E", x"EBCF", x"ECC4", x"EEB9",
		x"F288", x"F87D", x"0027", x"07F2", x"0E9C", x"12E1", x"147A", x"13C4",
		x"1182", x"0EC8", x"0C70", x"0ABE", x"0942", x"077E", x"04BB", x"00F3",
		x"FC53", x"F725", x"F232", x"EE3D", x"EC5D", x"ED3D", x"F108", x"F73F",
		x"FECD", x"06AD", x"0D74", x"1239", x"1462", x"13AD", x"105D", x"0AD8",
		x"03D2", x"FC51", x"F54A", x"EFD8", x"ECA9", x"EC48", x"EEB4", x"F36D",
		x"F9EB", x"012A", x"0865", x"0E73", x"1282", x"13FA", x"129D", x"0EC4",
		x"08B3", x"017C", x"F9E7", x"F32A", x"EE13", x"EB58", x"EB43", x"EDFB",
		x"F36E", x"FB0D", x"03A8", x"0B95", x"1120", x"134D", x"1218", x"0E80",
		x"0A09", x"0671", x"050B", x"0681", x"0A45", x"0EE9", x"1215", x"125D",
		x"0F38", x"08F7", x"0126", x"F937", x"F275", x"EDE6", x"EC22", x"ED07",
		x"F044", x"F57F", x"FC1E", x"037A", x"0A66", x"1004", x"135D", x"13F1",
		x"11DB", x"0D2A", x"0687", x"FED3", x"F765", x"F164", x"ED78", x"EBD9",
		x"ECD1", x"F07C", x"F6A0", x"FE77", x"06B7", x"0D99", x"11F1", x"12B4",
		x"0FFF", x"0B3B", x"0678", x"03CB", x"0484", x"0886", x"0DCC", x"11F8",
		x"12F9", x"10C0", x"0C5E", x"0814", x"058B", x"0621", x"0982", x"0E38",
		x"11C5", x"1234", x"0EF1", x"087D", x"007F", x"F854", x"F16B", x"ECCE",
		x"EAF0", x"EBE8", x"EF6F", x"F529", x"FC7D", x"04A5", x"0C03", x"1172",
		x"13F2", x"1341", x"1002", x"0B11", x"058E", x"002A", x"FB6E", x"F76B",
		x"F461", x"F20F", x"F048", x"EEF6", x"EE1C", x"ED4B", x"EC9F", x"EBEE",
		x"EB6D", x"EB25", x"EB17", x"EB7A", x"EC81", x"EEB0", x"F22A", x"F70D",
		x"FD29", x"0418", x"0AC8", x"1054", x"1380", x"1366", x"1016", x"0A30",
		x"02EE", x"FB8B", x"F4C4", x"EF9D", x"EC8D", x"EC19", x"EEC8", x"F490",
		x"FCB9", x"05C2", x"0D8C", x"125E", x"1421", x"1413", x"13B2", x"13AD",
		x"13C6", x"1292", x"0F19", x"0932", x"0148", x"F93A", x"F308", x"F0DE",
		x"F30F", x"F98C", x"0219", x"0A3C", x"1021", x"1349", x"1460", x"145F",
		x"1422", x"135A", x"1165", x"0D5A", x"06FC", x"FF13", x"F781", x"F283",
		x"F15C", x"F44F", x"FA4D", x"01F9", x"09BF", x"0FEC", x"1331", x"1348",
		x"10D7", x"0D45", x"0A01", x"075B", x"056A", x"03A8", x"0201", x"0028",
		x"FDFE", x"FBB4", x"F914", x"F650", x"F38F", x"F12C", x"EF5A", x"EE0A",
		x"ED29", x"EC5F", x"EBC6", x"EB47", x"EB1B", x"EB58", x"EBFD", x"ED03",
		x"EE70", x"F00B", x"F18D", x"F2EC", x"F42B", x"F57C", x"F73E", x"F9D3",
		x"FDAD", x"02D1", x"08E8", x"0E7A", x"1203", x"1232", x"0EE5", x"0966",
		x"03F6", x"0111", x"01D6", x"05E7", x"0B9F", x"10B0", x"130B", x"1207",
		x"0EB1", x"0ACC", x"0885", x"091E", x"0C33", x"102E", x"12C6", x"121B",
		x"0DA1", x"065C", x"FDE7", x"F600", x"EFEB", x"EC60", x"EB71", x"ED21",
		x"F0F8", x"F6EE", x"FE75", x"0695", x"0DBD", x"123F", x"1347", x"10CB",
		x"0C44", x"071C", x"02C8", x"0013", x"FF00", x"FF96", x"0143", x"0403",
		x"0734", x"0A80", x"0D10", x"0EB2", x"0FA1", x"0FB8", x"0EF3", x"0D09",
		x"0A19", x"0644", x"01B9", x"FCC0", x"F794", x"F2B4", x"EED2", x"ECA6",
		x"ECCC", x"EF96", x"F508", x"FC75", x"04B6", x"0C33", x"1187", x"13AC",
		x"12C4", x"0F6E", x"0A75", x"04AC", x"FEED", x"F9AD", x"F559", x"F1C2",
		x"EF2E", x"ED5B", x"EC77", x"EC2D", x"EC46", x"ECCD", x"EDD9", x"EFB4",
		x"F262", x"F569", x"F855", x"FA3E", x"FA5B", x"F833", x"F454", x"F016",
		x"ED6F", x"EE06", x"F241", x"F892", x"FE93", x"018F", x"0073", x"FB93",
		x"F4F3", x"EF7D", x"ED55", x"EEDC", x"F25E", x"F592", x"F66C", x"F470",
		x"F0D9", x"EDDA", x"EDD0", x"F1BB", x"F834", x"FEDF", x"03A6", x"0573",
		x"047D", x"019D", x"FDB9", x"F97B", x"F5C1", x"F2F3", x"F170", x"F186",
		x"F326", x"F5F1", x"F979", x"FD41", x"00BF", x"0368", x"04B9", x"049B",
		x"030B", x"004C", x"FCE4", x"F978", x"F672", x"F456", x"F2FC", x"F266",
		x"F2BC", x"F3D8", x"F5AA", x"F7F5", x"FACA", x"FDE4", x"0170", x"050C",
		x"0881", x"0BA7", x"0E4C", x"1062", x"11F9", x"1305", x"13A7", x"13C0",
		x"13A4", x"1342", x"1253", x"10B7", x"0E6B", x"0BEB", x"0986", x"07EA",
		x"0743", x"0779", x"08C3", x"0AC0", x"0D3D", x"0FB7", x"11D8", x"1350",
		x"1414", x"148F", x"14D7", x"14F3", x"14E8", x"14A8", x"13DD", x"124D",
		x"0F8B", x"0AF5", x"04B1", x"FD47", x"F600", x"F02B", x"ECCE", x"EC21",
		x"EDA3", x"F0ED", x"F4DD", x"F8B3", x"FBFD", x"FEB2", x"010E", x"02D8",
		x"0474", x"05BD", x"0705", x"08A8", x"0A87", x"0C9E", x"0EA4", x"10BF",
		x"12C0", x"142C", x"1496", x"136D", x"1074", x"0BD5", x"05BA", x"FE7C",
		x"F715", x"F0E9", x"ED73", x"EE03", x"F29B", x"F9ED", x"0243", x"09A5",
		x"0F10", x"123D", x"135D", x"1299", x"1000", x"0B9D", x"0552", x"FDA2",
		x"F607", x"F004", x"ED54", x"EED0", x"F42B", x"FC53", x"053B", x"0CCD",
		x"11E4", x"14A5", x"15DA", x"15DD", x"144F", x"10C8", x"0B08", x"036C",
		x"FB2B", x"F3A5", x"EE16", x"EB8D", x"EC41", x"EFC0", x"F590", x"FCFF",
		x"051D", x"0C94", x"1229", x"1525", x"15E9", x"1572", x"1500", x"14DF",
		x"14E4", x"1465", x"12C8", x"0FCE", x"0B3E", x"0535", x"FE2A", x"F713",
		x"F13A", x"ED6B", x"EC3C", x"ED8E", x"F07D", x"F474", x"F88C", x"FC0F",
		x"FEE0", x"012E", x"033F", x"0530", x"0728", x"0931", x"0B26", x"0D02",
		x"0EB1", x"1028", x"1199", x"12E8", x"1407", x"14A4", x"14D3", x"1453",
		x"1341", x"11E9", x"1073", x"0F77", x"0F21", x"0FB7", x"1129", x"131F",
		x"147E", x"13A9", x"0FAF", x"08CA", x"0053", x"F80C", x"F151", x"ECFC",
		x"EB45", x"EC31", x"EFAF", x"F557", x"FC99", x"0484", x"0BE1", x"10FC",
		x"127E", x"101F", x"0AA6", x"0405", x"FDBF", x"F94F", x"F7CD", x"F96A",
		x"FDDF", x"040D", x"0A8F", x"0FEC", x"1306", x"131F", x"1036", x"0B58",
		x"0594", x"0051", x"FC1D", x"F917", x"F74B", x"F6D0", x"F81D", x"FB89",
		x"0102", x"0795", x"0DDA", x"1210", x"134B", x"1204", x"0F7C", x"0D84",
		x"0D78", x"0F70", x"121F", x"1326", x"10BF", x"0AFB", x"031A", x"FB5A",
		x"F54F", x"F199", x"EFBE", x"EEEE", x"EEA7", x"EE1C", x"ED2C", x"EC08",
		x"EBB3", x"ED42", x"F1A7", x"F89A", x"00AA", x"0870", x"0EA0", x"12B1",
		x"14BC", x"1556", x"152B", x"14CC", x"142A", x"1323", x"115C", x"0EDD",
		x"0B8A", x"07CC", x"03CD", x"FF81", x"FB7B", x"F7F8", x"F59F", x"F4A0",
		x"F545", x"F7F5", x"FCF5", x"03D3", x"0AEA", x"1072", x"130D", x"12D8",
		x"1121", x"0FB3", x"0FBC", x"1137", x"12DD", x"12A9", x"0F42", x"08B8",
		x"009C", x"F8D1", x"F301", x"EF83", x"EDFF", x"ED76", x"ED20", x"EC8B",
		x"EB9E", x"EB17", x"EBA2", x"EE40", x"F346", x"FA7A", x"0281", x"09F4",
		x"0FC2", x"133F", x"14F9", x"1581", x"1566", x"14DC", x"13CF", x"1213",
		x"0FDA", x"0DBD", x"0C5D", x"0C4F", x"0D8E", x"0FC8", x"121A", x"13D4",
		x"14D3", x"155F", x"15AF", x"153D", x"1313", x"0E39", x"0725", x"FED7",
		x"F6FC", x"F0B4", x"EC93", x"EAC5", x"EB42", x"EDF5", x"F28F", x"F915",
		x"00EE", x"0904", x"0F87", x"1356", x"1466", x"13C2", x"1282", x"114F",
		x"102E", x"0F2F", x"0E16", x"0C86", x"0A96", x"081B", x"051E", x"01C2",
		x"FE4E", x"FB4C", x"F913", x"F7BB", x"F76C", x"F82C", x"F9F3", x"FCA3",
		x"0004", x"0373", x"0693", x"08D2", x"0A19", x"0A0F", x"0867", x"0551",
		x"0122", x"FCAC", x"F8DE", x"F688", x"F642", x"F895", x"FDB9", x"04CF",
		x"0C1B", x"113C", x"131B", x"11EE", x"0F97", x"0E47", x"0F00", x"1118",
		x"12E2", x"129C", x"0F18", x"08D2", x"016F", x"FB0A", x"F722", x"F5E7",
		x"F6F2", x"F979", x"FCFD", x"013C", x"057F", x"0958", x"0C7E", x"0EFA",
		x"10DC", x"1242", x"1322", x"139A", x"13F3", x"1457", x"1498", x"1483",
		x"13E3", x"12AA", x"110B", x"0F27", x"0D28", x"0B84", x"0ABE", x"0B0B",
		x"0C39", x"0E21", x"1027", x"1226", x"139B", x"149D", x"14E9", x"14FC",
		x"14A0", x"13BA", x"1210", x"0F81", x"0C8E", x"0A2C", x"0985", x"0AD5",
		x"0DBD", x"10ED", x"129B", x"1192", x"0D50", x"06EF", x"004B", x"FBEA",
		x"FB35", x"FE50", x"0444", x"0AFE", x"1046", x"1291", x"1183", x"0DCE",
		x"08D7", x"03D2", x"FFAE", x"FCD0", x"FAE5", x"F947", x"F79F", x"F5F2",
		x"F43A", x"F25E", x"F09B", x"EEE5", x"ED77", x"EC73", x"EBBE", x"EB4F",
		x"EB45", x"EB8F", x"EC39", x"ED40", x"EEEF", x"F128", x"F3A2", x"F5E2",
		x"F724", x"F6FE", x"F596", x"F373", x"F0F4", x"EEB6", x"ECE1", x"EB87",
		x"EAB2", x"EAFD", x"ED37", x"F211", x"F927", x"018E", x"0969", x"0F99",
		x"13C8", x"15EE", x"15FE", x"13DA", x"0F4E", x"0895", x"008C", x"F84F",
		x"F15D", x"ECDC", x"EB61", x"ECC3", x"F079", x"F627", x"FD9A", x"05E6",
		x"0D67", x"129B", x"14A2", x"1414", x"123C", x"106F", x"0F0E", x"0E09",
		x"0D33", x"0BE2", x"09F9", x"074B", x"03C4", x"FFE4", x"FBFD", x"F89D",
		x"F5E2", x"F445", x"F3AE", x"F40E", x"F535", x"F71B", x"F9CB", x"FCCC",
		x"FFD6", x"0257", x"0450", x"057A", x"05D5", x"055D", x"044E", x"02C6",
		x"00A7", x"FD93", x"F973", x"F49F", x"F00F", x"ED27", x"ED2B", x"F072",
		x"F65B", x"FD83", x"043F", x"08C8", x"0A19", x"07AB", x"01E8", x"FA9B",
		x"F3D3", x"EF2D", x"ED73", x"EE1C", x"EFE2", x"F1A6", x"F240", x"F159",
		x"EF5E", x"ED4C", x"EBDC", x"EB38", x"EB42", x"EBDA", x"ECB7", x"EDA7",
		x"EE71", x"EF39", x"F074", x"F2D2", x"F680", x"FBD0", x"026D", x"098D",
		x"0F92", x"131A", x"1371", x"110A", x"0D87", x"0A66", x"089F", x"086B",
		x"09DD", x"0C74", x"0F72", x"1231", x"1405", x"14FF", x"1525", x"149F",
		x"130C", x"1088", x"0D11", x"096B", x"06DA", x"0667", x"0875", x"0C52",
		x"106A", x"128A", x"115E", x"0CF5", x"069F", x"00D5", x"FE01", x"FF22",
		x"03F0", x"0A78", x"1016", x"12D3", x"1217", x"0EBC", x"0A99", x"0768",
		x"05E3", x"064D", x"0845", x"0B19", x"0E48", x"112E", x"137A", x"14D2",
		x"1549", x"1509", x"144E", x"136C", x"1268", x"1155", x"105F", x"0FC5",
		x"0FF2", x"10EC", x"127E", x"13E9", x"14F2", x"156B", x"156F", x"1546",
		x"151D", x"1521", x"151D", x"14BC", x"13D7", x"1252", x"10C6", x"0FC9",
		x"0FCA", x"10A7", x"1203", x"1366", x"1457", x"14D5", x"150B", x"154C",
		x"1598", x"152D", x"1344", x"0F13", x"0895", x"00B1", x"F8B4", x"F229",
		x"EDDF", x"EBCB", x"EB7E", x"EBFF", x"ED4E", x"EF50", x"F214", x"F55C",
		x"F8C9", x"FC27", x"FF38", x"01DE", x"0449", x"0670", x"089C", x"0AE2",
		x"0D2A", x"0F4C", x"1132", x"12C4", x"13F9", x"14AE", x"150A", x"152B",
		x"1535", x"14DE", x"13ED", x"1253", x"103C", x"0DD2", x"0B62", x"0972",
		x"0804", x"0714", x"06CF", x"06D6", x"0767", x"0848", x"09C7", x"0BE5",
		x"0EBD", x"11C3", x"141B", x"1473", x"11DE", x"0C83", x"054A", x"FD89",
		x"F6A5", x"F163", x"EE75", x"EE19", x"F020", x"F454", x"FA92", x"0225",
		x"0A01", x"1031", x"1307", x"11E8", x"0D21", x"0615", x"FE29", x"F6B7",
		x"F0DB", x"ED21", x"EBAA", x"EBFE", x"ED98", x"EFA7", x"F15D", x"F2B2",
		x"F3AF", x"F503", x"F708", x"FA87", x"FF99", x"061B", x"0C96", x"116F",
		x"1313", x"1155", x"0D2E", x"08A4", x"05C7", x"0547", x"0710", x"0A23",
		x"0D7A", x"104E", x"124B", x"130D", x"12B4", x"1110", x"0DDC", x"089A",
		x"0190", x"F987", x"F240", x"ED59", x"EC36", x"EF50", x"F5DF", x"FEC6",
		x"07A4", x"0EB6", x"12F9", x"14EE", x"1565", x"1559", x"150C", x"13B9",
		x"1083", x"0AF5", x"0344", x"FAC5", x"F342", x"EDFE", x"EB31", x"EA63",
		x"EABE", x"EB67", x"EC19", x"ECD8", x"ED81", x"EE55", x"EF55", x"F0A6",
		x"F233", x"F3DC", x"F5A1", x"F7C9", x"FAC0", x"FED0", x"042B", x"0A1D",
		x"0F5E", x"12B1", x"1309", x"1063", x"0B9D", x"062C", x"0195", x"FE9B",
		x"FD95", x"FE44", x"0034", x"0318", x"06BF", x"0B09", x"0F59", x"12A3",
		x"138A", x"113B", x"0BD6", x"0458", x"FC4B", x"F594", x"F1A2", x"F10F",
		x"F437", x"FA8B", x"0298", x"0A76", x"1065", x"13A9", x"14CD", x"14C0",
		x"1474", x"1426", x"12EF", x"0FAD", x"09D0", x"01DB", x"F99F", x"F330",
		x"EF4E", x"EDD1", x"EDEB", x"EF21", x"F16A", x"F4DD", x"F97F", x"FF28",
		x"052A", x"0AF1", x"0FB4", x"12AE", x"1375", x"11D0", x"0DC7", x"080E",
		x"01BC", x"FBE4", x"F703", x"F348", x"F0AD", x"EF0A", x"EE61", x"EE44",
		x"EE5C", x"EEC3", x"EF63", x"F044", x"F164", x"F2D8", x"F4C0", x"F74F",
		x"FAC6", x"FEFC", x"0363", x"0795", x"0B26", x"0DEA", x"0FC1", x"10BC",
		x"10BA", x"0FBE", x"0D78", x"0989", x"03E1", x"FCFA", x"F5D4", x"F010",
		x"ED01", x"ED9F", x"F1DF", x"F8BE", x"00A6", x"081B", x"0E37", x"1261",
		x"1483", x"1487", x"12AB", x"0F74", x"0B7A", x"075D", x"0398", x"00D9",
		x"FF76", x"000E", x"028B", x"0676", x"0B48", x"1006", x"1332", x"13A4",
		x"110C", x"0BEC", x"05A6", x"FF4F", x"F9A3", x"F4BB", x"F101", x"EE7E",
		x"ED0E", x"ECC1", x"ED6F", x"EFFB", x"F4E1", x"FC1B", x"0477", x"0C17",
		x"1176", x"1450", x"1542", x"154A", x"1534", x"1479", x"1284", x"0E64",
		x"07C5", x"FF77", x"F750", x"F128", x"ED9E", x"EC73", x"ECA8", x"EDE1",
		x"EFF5", x"F31F", x"F777", x"FCB5", x"0270", x"087F", x"0E0B", x"1241",
		x"1406", x"12DF", x"0F24", x"0996", x"037D", x"FDAA", x"F903", x"F5B4",
		x"F3B9", x"F292", x"F1C2", x"F0CB", x"EF7C", x"EE0D", x"EC92", x"EB85",
		x"EAEF", x"EAFD", x"EBC9", x"EC93", x"ECF9", x"ECBF", x"EC26", x"EB8F",
		x"EB4B", x"EB73", x"EBD6", x"EC56", x"ECA8", x"EC94", x"EC21", x"EBDD",
		x"ECB4", x"EFDC", x"F5B4", x"FDC8", x"0684", x"0DE9", x"12B7", x"1445",
		x"12EB", x"0F36", x"09E1", x"0344", x"FC21", x"F564", x"F01C", x"ED81",
		x"EE47", x"F245", x"F8C3", x"0013", x"06D7", x"0BFA", x"0F39", x"107D",
		x"1081", x"0F94", x"0DEE", x"0B90", x"0860", x"0494", x"0079", x"FC74",
		x"F876", x"F496", x"F12C", x"EE8F", x"ED0D", x"EC69", x"ECBF", x"EE91",
		x"F2B2", x"F979", x"01A0", x"0992", x"0FB2", x"1363", x"14FF", x"1577",
		x"1535", x"1452", x"1242", x"0E36", x"07EB", x"FFAB", x"F768", x"F0D0",
		x"ECD2", x"EB4E", x"EB82", x"EC7A", x"ED9C", x"EEA7", x"EEEC", x"EE47",
		x"ED0D", x"EC06", x"EC41", x"EEB1", x"F3CC", x"FB0D", x"0313", x"0A23",
		x"0EE1", x"10E8", x"10AD", x"0EE4", x"0BD7", x"0805", x"03D1", x"0019",
		x"FDD0", x"FD9B", x"FF71", x"02D6", x"071A", x"0B17", x"0E1A", x"0FEE",
		x"103C", x"0E9E", x"0A74", x"03D2", x"FBE8", x"F468", x"EF1E", x"EC71",
		x"EC32", x"ED32", x"EE6E", x"EF13", x"EEB8", x"ED9D", x"EC6A", x"EB9D",
		x"EB55", x"EBA9", x"ECCB", x"EE74", x"F056", x"F22E", x"F3D5", x"F594",
		x"F783", x"F9CF", x"FC59", x"FF82", x"02F5", x"069B", x"0A21", x"0CEE",
		x"0ED0", x"0FBB", x"0F98", x"0ED1", x"0D58", x"0AFD", x"0841", x"055A",
		x"0279", x"0032", x"FEDC", x"FE55", x"FE55", x"FECF", x"FFCF", x"018B",
		x"0452", x"083C", x"0CD7", x"1125", x"1396", x"1316", x"0F8B", x"09A7",
		x"0275", x"FB5E", x"F5E7", x"F34F", x"F44C", x"F86B", x"FEE4", x"0651",
		x"0D14", x"11DA", x"139A", x"1262", x"0F0B", x"0B2C", x"07AC", x"04F1",
		x"02BC", x"00F5", x"FF37", x"FD6B", x"FB99", x"F9AB", x"F7DE", x"F608",
		x"F420", x"F224", x"EFFC", x"EDB7", x"EBFF", x"EBA2", x"ED9F", x"F25B",
		x"F969", x"015E", x"08D4", x"0EA7", x"1266", x"141D", x"141A", x"12C1",
		x"1033", x"0CD0", x"093D", x"067C", x"058E", x"0729", x"0AD2", x"0F2E",
		x"120D", x"11A6", x"0D88", x"0745", x"0169", x"FE7C", x"FFEB", x"050F",
		x"0BA6", x"10B9", x"1283", x"10C5", x"0D48", x"0A65", x"09CF", x"0BE0",
		x"0F86", x"123D", x"1240", x"0EB9", x"08F9", x"02C2", x"FDD8", x"FB3F",
		x"FB0A", x"FCE4", x"0029", x"041C", x"0812", x"0BB9", x"0EAA", x"10F8",
		x"129A", x"139C", x"1453", x"14BA", x"14D9", x"14DD", x"148B", x"13D2",
		x"1273", x"10B2", x"0E94", x"0C51", x"0A44", x"0892", x"0794", x"0748",
		x"07ED", x"095A", x"0B20", x"0CF3", x"0EB5", x"108E", x"1258", x"13D7",
		x"14D1", x"14D3", x"13F6", x"127B", x"10E4", x"0FA4", x"0F81", x"1077",
		x"1208", x"1339", x"12E8", x"1020", x"0AC3", x"03B3", x"FC71", x"F6FE",
		x"F4D6", x"F661", x"FB53", x"0262", x"09A8", x"0F7E", x"126D", x"1223",
		x"0F51", x"0B57", x"07A5", x"0535", x"040F", x"0322", x"01D4", x"FF46",
		x"FB51", x"F682", x"F1BF", x"EE2B", x"ED00", x"EEA3", x"F2CB", x"F87F",
		x"FEF9", x"0505", x"0A2C", x"0E07", x"10D4", x"12BC", x"13E8", x"1480",
		x"14DA", x"14C2", x"141A", x"12F1", x"1113", x"0E74", x"0B90", x"0916",
		x"07D3", x"088E", x"0B25", x"0ED3", x"11F4", x"1330", x"111F", x"0C06",
		x"0593", x"000E", x"FD93", x"FEBF", x"0302", x"08DE", x"0E71", x"1215",
		x"126F", x"0F00", x"085B", x"FFDB", x"F7A2", x"F121", x"ED30", x"EBDC",
		x"ECDC", x"EFD5", x"F446", x"F970", x"FE7E", x"02CB", x"0627", x"08CB",
		x"0AEC", x"0C65", x"0D0D", x"0C93", x"0AC8", x"0818", x"050C", x"01D3",
		x"FEA5", x"FBE8", x"FA1A", x"F99E", x"FA91", x"FCDD", x"0011", x"03B6",
		x"0746", x"09F2", x"0B64", x"0B53", x"097B", x"05AB", x"FFFC", x"F938",
		x"F299", x"EDF1", x"EC7F", x"EEE9", x"F4DD", x"FCFB", x"0576", x"0CD3",
		x"11C4", x"13F6", x"13AD", x"11FA", x"1026", x"0F17", x"0F31", x"1051",
		x"11FC", x"13AC", x"14C4", x"1544", x"155E", x"157C", x"1594", x"1577",
		x"14F7", x"1408", x"12AA", x"1105", x"0ED2", x"0BF9", x"0882", x"048C",
		x"00A1", x"FD0F", x"FA2A", x"F852", x"F81A", x"F9D6", x"FE05", x"03F6",
		x"0A99", x"1021", x"1313", x"12BC", x"1002", x"0C91", x"09EE", x"0938",
		x"0A58", x"0CF6", x"0FFA", x"128C", x"1451", x"150F", x"151D", x"14A0",
		x"1396", x"11E6", x"0F78", x"0CB5", x"0A8F", x"09EB", x"0B42", x"0DFC",
		x"1116", x"1356", x"1357", x"108D", x"0B02", x"03E0", x"FC88", x"F65A",
		x"F1B4", x"EE92", x"ECBD", x"EBE2", x"EBA9", x"EB7E", x"EB4D", x"EB0D",
		x"EB26", x"EB95", x"EC5A", x"ED37", x"EE34", x"EFEA", x"F258", x"F582",
		x"F8F6", x"FC69", x"FFC4", x"032B", x"0657", x"08E0", x"0A4C", x"0AB8",
		x"0A0F", x"080F", x"050B", x"0146", x"FD97", x"FA8B", x"F895", x"F81B",
		x"F9C6", x"FDD1", x"03CD", x"0A59", x"0FE9", x"1338", x"13B1", x"1136",
		x"0CB4", x"0719", x"0154", x"FC54", x"F878", x"F5F4", x"F4C6", x"F4EC",
		x"F675", x"F99E", x"FE7F", x"04AC", x"0B17", x"1051", x"131C", x"12EE",
		x"0FEE", x"0B42", x"0666", x"0286", x"FFD7", x"FE0B", x"FCB1", x"FB3D",
		x"F95C", x"F72D", x"F4A5", x"F1EE", x"EF48", x"ED2D", x"EBB9", x"EAF2",
		x"EA7D", x"EA80", x"EB68", x"EE24", x"F2E8", x"F9A0", x"0182", x"0959",
		x"0FBA", x"13D4", x"1548", x"150C", x"1422", x"1341", x"1274", x"1176",
		x"0FEC", x"0D83", x"09FF", x"04FF", x"FEFE", x"F85C", x"F243", x"EDBB",
		x"EBE4", x"ED44", x"F202", x"F956", x"01D5", x"0A0D", x"1048", x"1395",
		x"13D6", x"11FE", x"0F9F", x"0DB5", x"0D2C", x"0E15", x"0FE9", x"1209",
		x"13C1", x"14CE", x"1544", x"1539", x"1481", x"129D", x"0EC8", x"08A7",
		x"00AE", x"F82F", x"F0F9", x"ECCC", x"EC5B", x"EF21", x"F431", x"FA86",
		x"0146", x"080C", x"0DF4", x"124B", x"13F7", x"1224", x"0CC6", x"0503",
		x"FC8C", x"F51C", x"EFCA", x"ECAF", x"EB5E", x"EB05", x"EB47", x"EBC5",
		x"ECE1", x"EE93", x"F0C1", x"F2F7", x"F4B4", x"F59B", x"F5BD", x"F509",
		x"F398", x"F1A6", x"EFA6", x"ED98", x"EC19", x"EBF0", x"EE06", x"F318",
		x"FA69", x"02A8", x"09EA", x"0F7D", x"12F9", x"1483", x"1409", x"118D",
		x"0CDE", x"0634", x"FE42", x"F643", x"EFE0", x"EC33", x"EB58", x"EC8D",
		x"EEA4", x"F0EF", x"F2E2", x"F446", x"F510", x"F528", x"F499", x"F357",
		x"F171", x"EF43", x"ED75", x"EC14", x"EB37", x"EAA0", x"EAAC", x"EC48",
		x"F03C", x"F673", x"FE61", x"06AD", x"0DC0", x"129F", x"150D", x"15A8",
		x"1550", x"14A1", x"1396", x"1215", x"0FFD", x"0E1B", x"0D68", x"0E60",
		x"10B2", x"12CB", x"1310", x"1003", x"09F3", x"023E", x"FAD9", x"F5CD",
		x"F3A9", x"F410", x"F643", x"F9B5", x"FDBF", x"01D4", x"0547", x"0768",
		x"07A5", x"0646", x"03B2", x"0090", x"FD2C", x"F9AF", x"F6C5", x"F4BF",
		x"F3DC", x"F42D", x"F59D", x"F7E0", x"FAD8", x"FE1A", x"01A3", x"04FB",
		x"07F3", x"0A55", x"0C68", x"0E44", x"100D", x"11AF", x"1307", x"1414",
		x"14C9", x"153B", x"1542", x"14E1", x"144C", x"137F", x"1294", x"1161",
		x"0F9D", x"0D51", x"0A90", x"07AF", x"0499", x"01A8", x"FEE9", x"FCB9",
		x"FB13", x"FA02", x"F9B4", x"FA2A", x"FB90", x"FDE8", x"013B", x"04EB",
		x"089B", x"0C49", x"0FC7", x"1290", x"13C6", x"1299", x"0EB7", x"08A2",
		x"012F", x"F965", x"F284", x"EDAF", x"EBE3", x"ED10", x"F0BF", x"F662",
		x"FD48", x"04D3", x"0BD5", x"1107", x"136E", x"12E7", x"0F90", x"09C9",
		x"02B3", x"FB86", x"F593", x"F153", x"EEC2", x"ED3E", x"EC52", x"EBE5",
		x"EB6E", x"EAE6", x"EA9C", x"EBEF", x"EFE7", x"F6C1", x"FF77", x"07E5",
		x"0E88", x"12C9", x"1513", x"15E3", x"154C", x"12D9", x"0E35", x"0776",
		x"FF46", x"F716", x"F0A5", x"ECEB", x"EBD6", x"ED52", x"F0E5", x"F6B1",
		x"FE32", x"066F", x"0D9A", x"1200", x"1229", x"0DED", x"066C", x"FDB8",
		x"F5E1", x"EFFA", x"EC69", x"EAA0", x"EA2C", x"EAA0", x"EC14", x"EEFA",
		x"F449", x"FBBF", x"046B", x"0C34", x"11C0", x"145E", x"14F6", x"1450",
		x"1337", x"123C", x"1188", x"10FC", x"10AB", x"10A1", x"10A7", x"10D2",
		x"1126", x"11F4", x"1338", x"1478", x"1510", x"141E", x"110C", x"0BF7",
		x"0522", x"FD57", x"F5DE", x"F009", x"EC81", x"EB5F", x"EBF6", x"ED79",
		x"EF22", x"F084", x"F1AC", x"F2C0", x"F4A4", x"F7C1", x"FC60", x"0293",
		x"0981", x"0F8A", x"130B", x"1303", x"0FCB", x"0B60", x"07D8", x"06A5",
		x"07E5", x"0AE8", x"0E4A", x"1120", x"1306", x"141D", x"1412", x"125E",
		x"0E1D", x"073D", x"FED8", x"F6BF", x"F090", x"ECC0", x"EAF1", x"EA68",
		x"EAAB", x"EBFE", x"EEF5", x"F43A", x"FBDB", x"04B0", x"0CBF", x"1215",
		x"13C4", x"11C3", x"0CBE", x"0610", x"FEC8", x"F7DC", x"F241", x"EE40",
		x"EBD3", x"EACD", x"EAC3", x"EB27", x"EBCC", x"ECB5", x"ED9F", x"EEA2",
		x"EFF0", x"F17B", x"F33B", x"F56B", x"F7B3", x"FA0C", x"FCAF", x"FF87",
		x"02BB", x"0652", x"09F0", x"0D3C", x"1003", x"1203", x"1329", x"138B",
		x"130F", x"1184", x"0EAF", x"0A05", x"0391", x"FC09", x"F4CB", x"EF41",
		x"ECB8", x"EE2A", x"F39C", x"FBE1", x"04DE", x"0CA4", x"11D8", x"14A0",
		x"157C", x"156C", x"14CF", x"1313", x"0F79", x"097F", x"01B0", x"F958",
		x"F25B", x"EE22", x"ED39", x"EFA0", x"F482", x"FB4B", x"032A", x"0AC8",
		x"1091", x"1352", x"12E4", x"1050", x"0CC0", x"092B", x"0628", x"0408",
		x"02F7", x"03B5", x"0629", x"0A03", x"0E69", x"11FB", x"1385", x"121B",
		x"0DE4", x"0807", x"0275", x"FE7A", x"FCF3", x"FDB9", x"0058", x"03EF",
		x"0804", x"0BEE", x"0F46", x"11AC", x"1304", x"1390", x"13CB", x"1421",
		x"149D", x"1506", x"14A9", x"12EE", x"0F1F", x"092D", x"0185", x"F957",
		x"F25B", x"EDA6", x"EB5F", x"EB14", x"EBAA", x"EC44", x"EC6F", x"EC0E",
		x"EB8D", x"EB72", x"EC2B", x"EDA8", x"EF93", x"F16A", x"F30A", x"F445",
		x"F559", x"F6A6", x"F8CF", x"FC7E", x"01BD", x"07D7", x"0DC1", x"119B",
		x"1235", x"0F70", x"0A78", x"059A", x"02E0", x"034B", x"06A7", x"0BA3",
		x"1056", x"12BA", x"11EB", x"0E33", x"0937", x"0499", x"018C", x"008C",
		x"018C", x"0423", x"0792", x"0B96", x"0F97", x"12D4", x"1415", x"1296",
		x"0DFD", x"0716", x"FF64", x"F829", x"F280", x"EF2B", x"EED8", x"F1EA",
		x"F7F3", x"FFB3", x"078C", x"0E35", x"12C4", x"14C2", x"149E", x"13A2",
		x"1318", x"1393", x"1448", x"1481", x"13EB", x"1311", x"1280", x"128F",
		x"1332", x"13F3", x"146B", x"1450", x"13E8", x"13A9", x"13B5", x"13F4",
		x"13CE", x"1267", x"0EF9", x"0902", x"0137", x"F90E", x"F273", x"EE0E",
		x"EBF4", x"EB4B", x"EB72", x"EBED", x"EC7F", x"ECD9", x"ECED", x"ECE1",
		x"ECB5", x"EC16", x"EB54", x"EACA", x"EACB", x"EB61", x"EC53", x"ED00",
		x"ED0F", x"ECA3", x"EC12", x"EB86", x"EB41", x"EB84", x"EC1F", x"ECDE",
		x"ED32", x"ECCA", x"EBDF", x"EB20", x"EAED", x"EB7B", x"EC4D", x"EC79",
		x"EC08", x"EB4C", x"EB6C", x"ED42", x"F19F", x"F85F", x"0094", x"08AE",
		x"0F11", x"1306", x"14E0", x"1563", x"1547", x"14D3", x"142E", x"13AB",
		x"134F", x"134B", x"1380", x"13EE", x"145F", x"14BF", x"14FF", x"14B2",
		x"13E7", x"128A", x"10C1", x"0ED0", x"0CD6", x"0B0A", x"093F", x"0766",
		x"0530", x"025B", x"FEDE", x"FAC3", x"F6B9", x"F333", x"F065", x"EE7B",
		x"EDAA", x"EDDE", x"EF77", x"F2CD", x"F847", x"FF78", x"071B", x"0DDD",
		x"126D", x"140F", x"12F4", x"1007", x"0C3F", x"086A", x"0500", x"02AD",
		x"0176", x"01AD", x"033E", x"05F9", x"09BB", x"0DE2", x"1193", x"1335",
		x"11CF", x"0D39", x"063C", x"FE08", x"F631", x"F024", x"ECAC", x"EC0D",
		x"EE1A", x"F20D", x"F74B", x"FD4D", x"034C", x"08A1", x"0CF1", x"0FD8",
		x"118B", x"1288", x"12E8", x"124A", x"101E", x"0BD3", x"057D", x"FE12",
		x"F6C5", x"F0CE", x"ED1C", x"EC16", x"ED4C", x"EF80", x"F18B", x"F2CE",
		x"F3A8", x"F4A4", x"F688", x"F99F", x"FE72", x"0486", x"0AFA", x"103B",
		x"12AA", x"11C5", x"0E31", x"09F9", x"072E", x"0709", x"09B9", x"0DD0",
		x"1168", x"1289", x"1077", x"0BCE", x"063B", x"0149", x"FE0C", x"FD07",
		x"FE40", x"0145", x"058D", x"0A76", x"0F0E", x"1297", x"146A", x"1481",
		x"12AD", x"0F1D", x"098F", x"025C", x"FA65", x"F325", x"EE3C", x"EC76",
		x"EE0E", x"F25E", x"F891", x"FF6C", x"05F8", x"0BA1", x"0FF5", x"130D",
		x"14B5", x"1541", x"152F", x"14BA", x"1424", x"1398", x"1369", x"139F",
		x"141B", x"1475", x"1442", x"135C", x"1272", x"121E", x"12A3", x"1394",
		x"1467", x"1441", x"1274", x"0E70", x"07E2", x"FF84", x"F6FA", x"F04C",
		x"ED34", x"EE53", x"F31D", x"F9EF", x"0131", x"0773", x"0BDF", x"0D9A",
		x"0C21", x"0798", x"00B0", x"F8EE", x"F279", x"EE4C", x"ECB3", x"ECF9",
		x"EDF1", x"EE7B", x"EE0B", x"ECDA", x"EB79", x"EAF6", x"EB0E", x"EB6D",
		x"EBCD", x"EBC6", x"EB8E", x"EB8F", x"EC37", x"ED47", x"EE3F", x"EE78",
		x"EDCB", x"ECE2", x"ECA0", x"EE1D", x"F1E2", x"F816", x"FFAD", x"070C",
		x"0C59", x"0F38", x"1017", x"0F67", x"0DB8", x"0AFB", x"075C", x"0347",
		x"FF30", x"FB4F", x"F7D5", x"F4C9", x"F222", x"EFFE", x"EE58", x"ED32",
		x"EC82", x"EC3F", x"ECAB", x"EDBE", x"EF4E", x"F142", x"F398", x"F63C",
		x"F8B9", x"FA65", x"FAAC", x"F98C", x"F75C", x"F4BB", x"F20B", x"EFA1",
		x"EDDA", x"EC90", x"EC0D", x"EBF8", x"EC36", x"ECD7", x"EE04", x"EFE9",
		x"F2E1", x"F6F3", x"FC0E", x"024B", x"090C", x"0F15", x"12E6", x"1387",
		x"1162", x"0D80", x"0968", x"0675", x"0566", x"064B", x"0874", x"0B3C",
		x"0E18", x"10A1", x"12C0", x"1423", x"14CB", x"14E7", x"14CE", x"145E",
		x"1390", x"126F", x"1108", x"0F86", x"0DDC", x"0C39", x"0ACD", x"0968",
		x"07E9", x"0595", x"01ED", x"FCF4", x"F73F", x"F1D5", x"EDED", x"ECAB",
		x"EE4B", x"F288", x"F802", x"FD41", x"015A", x"03D6", x"04CF", x"0462",
		x"02B4", x"FFB3", x"FB7A", x"F691", x"F1A5", x"EE39", x"ED20", x"EEF5",
		x"F387", x"F9D9", x"0070", x"061F", x"09E5", x"0AC3", x"08D6", x"040B",
		x"FD68", x"F660", x"F078", x"ED79", x"EE6C", x"F393", x"FB58", x"03E4",
		x"0B5A", x"10B6", x"1396", x"144E", x"1377", x"11CF", x"1044", x"0F23",
		x"0F0E", x"0FF7", x"117D", x"131B", x"140D", x"13B2", x"1190", x"0D87",
		x"07AB", x"008B", x"F94A", x"F2F1", x"EE3C", x"EBB7", x"EB81", x"ED3E",
		x"F03F", x"F3BC", x"F6C9", x"F8F5", x"F990", x"F89E", x"F643", x"F314",
		x"EF8E", x"ECB8", x"EBF1", x"EDD9", x"F279", x"F910", x"0020", x"06AC",
		x"0BF7", x"0FF6", x"129E", x"1415", x"1485", x"1455", x"13E5", x"12C8",
		x"10A0", x"0CBD", x"0735", x"0062", x"F906", x"F242", x"ED96", x"EC62",
		x"EEF3", x"F4B6", x"FC60", x"0480", x"0B9E", x"10E1", x"13F0", x"1521",
		x"14EF", x"13C9", x"121C", x"10AD", x"0F66", x"0E23", x"0C2F", x"0914",
		x"049E", x"FECD", x"F843", x"F253", x"EE33", x"ECC1", x"EE45", x"F201",
		x"F6EE", x"FBAC", x"FF6E", x"01A0", x"02B6", x"037A", x"04E7", x"07C3",
		x"0BAA", x"0F99", x"122F", x"1232", x"0F21", x"0981", x"0255", x"FB69",
		x"F6CF", x"F5D6", x"F90F", x"FF83", x"0753", x"0E17", x"1224", x"1337",
		x"1235", x"10CF", x"1062", x"114D", x"129F", x"1275", x"0EF8", x"0840",
		x"FF81", x"F70B", x"F05C", x"EC73", x"EB6F", x"ED50", x"F17A", x"F787",
		x"FEBD", x"063E", x"0D16", x"1206", x"140E", x"12E1", x"0EE7", x"08EE",
		x"022F", x"FB8B", x"F5F1", x"F1AF", x"EEC3", x"ECD6", x"EB7C", x"EABB",
		x"EA55", x"EA54", x"EA87", x"EACD", x"EAFB", x"EB0E", x"EB1E", x"EB92",
		x"EC9F", x"EE82", x"F147", x"F561", x"FACD", x"0147", x"0828", x"0E1E",
		x"1220", x"1375", x"1194", x"0D04", x"0670", x"FEE9", x"F786", x"F181",
		x"ED63", x"EBD8", x"ECF7", x"F0BF", x"F716", x"FF2D", x"0797", x"0E82",
		x"12C2", x"13D1", x"12A2", x"107C", x"0E9C", x"0DF5", x"0EDA", x"10B4",
		x"12B4", x"1442", x"1527", x"159F", x"15A4", x"1461", x"10D4", x"0AC8",
		x"02C7", x"FA53", x"F2DD", x"ED55", x"EA58", x"EA6A", x"ED9E", x"F398",
		x"FB73", x"03C6", x"0B4A", x"1104", x"1477", x"15BD", x"1517", x"1283",
		x"0DE1", x"06E7", x"FE66", x"F5CD", x"EF2A", x"EBAD", x"EB06", x"EC38",
		x"EDF4", x"EF77", x"F098", x"F154", x"F1D8", x"F23D", x"F268", x"F201",
		x"F0DE", x"EF4D", x"EDE7", x"ECB5", x"EBB7", x"EB45", x"EB3B", x"EBE1",
		x"ECE8", x"EE21", x"EF5C", x"F0A3", x"F1FE", x"F32A", x"F403", x"F43B",
		x"F3CF", x"F2E6", x"F195", x"EFDC", x"EDE0", x"EBFD", x"EB08", x"EBE1",
		x"EF22", x"F503", x"FCB2", x"04D6", x"0BDB", x"10E3", x"13CD", x"14FA",
		x"152C", x"14C4", x"13EE", x"1264", x"1014", x"0D8F", x"0BE1", x"0BEC",
		x"0DCF", x"10AC", x"12E5", x"12BF", x"0F68", x"0920", x"0184", x"FA5D",
		x"F4C5", x"F149", x"EF68", x"EE81", x"EDFE", x"ED6A", x"EC95", x"EBCE",
		x"EBED", x"EDEC", x"F264", x"F947", x"013A", x"08E4", x"0EEA", x"12BB",
		x"149F", x"150E", x"14F5", x"14B2", x"141A", x"12E9", x"10E8", x"0E42",
		x"0B8D", x"0924", x"070A", x"0520", x"033A", x"010E", x"FE81", x"FB99",
		x"F803", x"F410", x"F029", x"ED23", x"EBF4", x"ED19", x"F11F", x"F798",
		x"FF90", x"0795", x"0E30", x"126B", x"13B5", x"1202", x"0D8F", x"076E",
		x"00CE", x"FA9F", x"F5B7", x"F261", x"F03D", x"EEE4", x"EDD4", x"ECEC",
		x"EBE3", x"EB02", x"EB37", x"ED7C", x"F28C", x"FA1C", x"0282", x"0A3F",
		x"1075", x"148A", x"1615", x"149A", x"1042", x"0997", x"01A8", x"F968",
		x"F20A", x"ECA0", x"E9CE", x"E9E7", x"ECBC", x"F201", x"F956", x"01C3",
		x"09CE", x"109B", x"14DE", x"1615", x"1401", x"0EC0", x"0779", x"FF38",
		x"F754", x"F0C9", x"EC58", x"EA3A", x"EA67", x"EC9A", x"F0C0", x"F6D7",
		x"FEA6", x"0710", x"0E44", x"12F7", x"14B4", x"1452", x"12E9", x"114B",
		x"0FD0", x"0EA4", x"0DFB", x"0DB4", x"0DC1", x"0E22", x"0EE6", x"1043",
		x"11CB", x"131D", x"1412", x"1499", x"14D1", x"14A1", x"13F1", x"12C2",
		x"1159", x"0FAF", x"0DD3", x"0BC4", x"09A5", x"075B", x"0555", x"0353",
		x"0182", x"FF89", x"FD4F", x"FA41", x"F664", x"F21B", x"EE7C", x"ECAF",
		x"EDB3", x"F1B6", x"F80E", x"FF7E", x"05EB", x"09F6", x"0B3D", x"0A5C",
		x"07E2", x"047C", x"00A7", x"FCF1", x"FA55", x"F99B", x"FB5A", x"FF88",
		x"054B", x"0B70", x"1064", x"12B0", x"117A", x"0CFD", x"0634", x"FE4D",
		x"F6F4", x"F118", x"ED48", x"EBD0", x"ECC9", x"F065", x"F673", x"FE36",
		x"068B", x"0DC5", x"1284", x"1402", x"12AF", x"0FB4", x"0C7C", x"0A28",
		x"0916", x"099E", x"0B67", x"0DE1", x"1078", x"12B9", x"1450", x"1520",
		x"152F", x"14E1", x"1499", x"147A", x"143F", x"1358", x"112A", x"0D40",
		x"0735", x"FF60", x"F71E", x"F04D", x"EC81", x"EBC5", x"ECC9", x"EE06",
		x"EE28", x"ED52", x"EC68", x"ECE3", x"EFFC", x"F5DE", x"FD95", x"0599",
		x"0C53", x"1115", x"13B7", x"14AE", x"14A5", x"1465", x"146D", x"14CE",
		x"1520", x"141C", x"1102", x"0B92", x"045C", x"FC59", x"F4E2", x"EEFB",
		x"EB9A", x"EB4B", x"EE0E", x"F3AB", x"FB37", x"03BD", x"0BB1", x"118C",
		x"14BD", x"15A5", x"154F", x"14CD", x"1450", x"134B", x"11BF", x"0FDD",
		x"0EFF", x"0FAC", x"116C", x"12EF", x"1295", x"0FA2", x"09F7", x"02E3",
		x"FBCA", x"F646", x"F306", x"F204", x"F293", x"F466", x"F724", x"FAA1",
		x"FE94", x"02BD", x"069D", x"0A25", x"0D37", x"0FBE", x"11A4", x"12DE",
		x"13A0", x"1404", x"1404", x"139D", x"12C4", x"118F", x"0FF9", x"0DE8",
		x"0BAE", x"09A2", x"0819", x"074B", x"0785", x"08F2", x"0B54", x"0E0C",
		x"107D", x"1247", x"1362", x"1432", x"14C4", x"1538", x"1570", x"1550",
		x"14BB", x"1392", x"119A", x"0E30", x"08DB", x"01BD", x"F9E1", x"F2EB",
		x"EE37", x"EC43", x"EC98", x"EDEE", x"EF42", x"EFDA", x"EF79", x"EE56",
		x"ECE2", x"EBA5", x"EAFA", x"EB2F", x"EBDA", x"ECD3", x"EDCC", x"EE9A",
		x"EFA7", x"F158", x"F401", x"F790", x"FC02", x"0156", x"0732", x"0CFE",
		x"118D", x"13F1", x"134A", x"0F7C", x"08D4", x"00B7", x"F88C", x"F1D1",
		x"ED74", x"EC1D", x"ED9A", x"F0EA", x"F4D3", x"F7F0", x"F9C5", x"FA2F",
		x"F9A0", x"F815", x"F5BB", x"F2A0", x"EF4F", x"EC8A", x"EBE9", x"EE60",
		x"F3F6", x"FBBC", x"0401", x"0B50", x"10AB", x"1359", x"12BD", x"0EE1",
		x"0838", x"002C", x"F81F", x"F190", x"ECF4", x"EA60", x"E9A3", x"EA77",
		x"ECD0", x"F139", x"F7E8", x"0026", x"08A8", x"0F89", x"138D", x"1494",
		x"1387", x"1150", x"0E7B", x"0B45", x"082C", x"0637", x"0621", x"0840",
		x"0BF3", x"0FFD", x"12C3", x"1308", x"1026", x"0AA9", x"03C2", x"FD11",
		x"F78A", x"F363", x"F092", x"EECF", x"EDB5", x"ED3E", x"ED03", x"ED05",
		x"ED30", x"EDC6", x"EED5", x"F03C", x"F229", x"F4AD", x"F7B3", x"FB3D",
		x"FEA3", x"01B3", x"0495", x"074C", x"09D3", x"0BF2", x"0D91", x"0E88",
		x"0EFE", x"0EFB", x"0EAD", x"0DD9", x"0C5D", x"0A0C", x"06C7", x"0237",
		x"FCA7", x"F698", x"F109", x"ED12", x"EB7E", x"ECAF", x"F08A", x"F649",
		x"FCC1", x"031B", x"0887", x"0CCC", x"0FCB", x"11CE", x"131F", x"13B1",
		x"1357", x"11C8", x"0E7E", x"0940", x"0255", x"FAA9", x"F376", x"EE64",
		x"EC09", x"EC2C", x"EDE9", x"EFFE", x"F1AF", x"F2D4", x"F3E1", x"F564",
		x"F7CC", x"FBBB", x"0122", x"0774", x"0D7E", x"1173", x"1233", x"0FDA",
		x"0BB1", x"07F4", x"067E", x"083D", x"0C38", x"1095", x"12F5", x"11E7",
		x"0D74", x"0717", x"007D", x"FAE4", x"F6E3", x"F46B", x"F30C", x"F215",
		x"F0F8", x"EF5B", x"ED67", x"EBC6", x"EB4D", x"ECC8", x"F09F", x"F6B1",
		x"FE5D", x"065E", x"0D4D", x"11EC", x"135B", x"11A6", x"0D4F", x"073E",
		x"0070", x"F9C9", x"F3E7", x"EF64", x"EC8C", x"EB6B", x"EB8E", x"EC8D",
		x"EDE4", x"EEED", x"EED7", x"ED91", x"EC09", x"EBA7", x"EDF4", x"F2EC",
		x"F9F5", x"0194", x"0875", x"0D40", x"0F35", x"0E21", x"0A38", x"0419",
		x"FC9F", x"F52F", x"EF6D", x"ECFA", x"EEF3", x"F4C8", x"FD2E", x"0617",
		x"0DA8", x"127C", x"1483", x"14A3", x"1427", x"13D8", x"13BA", x"12B1",
		x"0F8E", x"09DB", x"026C", x"FA84", x"F3D3", x"EF71", x"ED7C", x"ED82",
		x"EEE5", x"F13B", x"F451", x"F804", x"FC28", x"002B", x"0423", x"07E6",
		x"0B58", x"0E12", x"102C", x"117F", x"122E", x"11C3", x"0FDF", x"0BC5",
		x"05A2", x"FE6E", x"F755", x"F16A", x"EDAC", x"ECA9", x"EDF4", x"F0AE",
		x"F394", x"F5DA", x"F751", x"F85C", x"F993", x"FB65", x"FE08", x"0178",
		x"0573", x"096D", x"0D06", x"0FA8", x"1155", x"11F5", x"1163", x"0F1E",
		x"0A44", x"0328", x"FB09", x"F39F", x"EE74", x"EC20", x"EBC1", x"EC4E",
		x"ECB9", x"EC73", x"EBBB", x"EB2D", x"EB20", x"EB9D", x"EC0C", x"EC08",
		x"EB7A", x"EB1C", x"EC0B", x"EF49", x"F53F", x"FD66", x"0647", x"0DD2",
		x"1286", x"13A4", x"1117", x"0B88", x"0418", x"FC89", x"F628", x"F1CF",
		x"EF80", x"EED0", x"EF42", x"F0D4", x"F359", x"F6B9", x"FA21", x"FD18",
		x"FF0D", x"FF9A", x"FED6", x"FCBC", x"F9CA", x"F687", x"F361", x"F096",
		x"EEA2", x"ED27", x"EC38", x"EB88", x"EB1E", x"EAD6", x"EAC8", x"EB2A",
		x"EC42", x"EEEE", x"F374", x"FA0D", x"01EB", x"09AE", x"0FC9", x"1368",
		x"14A9", x"14A0", x"1430", x"1420", x"1475", x"14CC", x"148A", x"13BA",
		x"12B6", x"1205", x"122B", x"12EC", x"13E6", x"14B7", x"14EE", x"148F",
		x"13ED", x"13BE", x"1422", x"147C", x"13D6", x"1177", x"0CB9", x"05B9",
		x"FD76", x"F564", x"EF25", x"EC43", x"ED61", x"F201", x"F8D1", x"003A",
		x"06EA", x"0C3B", x"0FF4", x"1213", x"12AE", x"123F", x"10EF", x"0EE6",
		x"0C29", x"08EA", x"0561", x"01CD", x"FE16", x"FA88", x"F754", x"F46B",
		x"F21A", x"F091", x"EFCA", x"EFA9", x"F04E", x"F21E", x"F4F0", x"F86D",
		x"FC02", x"FEE2", x"008E", x"004B", x"FDB5", x"F90C", x"F372", x"EEAD",
		x"ECA0", x"EE40", x"F283", x"F791", x"FB2C", x"FC31", x"FA9E", x"F72A",
		x"F34C", x"F01D", x"EDF1", x"ED02", x"ED8B", x"F012", x"F4D1", x"FBB0",
		x"03B8", x"0B4A", x"110C", x"1443", x"153B", x"14D8", x"1442", x"1407",
		x"1437", x"1460", x"143F", x"1387", x"1233", x"1053", x"0DF3", x"0B15",
		x"083B", x"055F", x"02CB", x"00C0", x"FF47", x"FE90", x"FEA9", x"FFBC",
		x"018F", x"0405", x"06C5", x"09A2", x"0C69", x"0EE2", x"10D4", x"1248",
		x"1354", x"143F", x"14CF", x"1510", x"14DB", x"1456", x"137F", x"129E",
		x"1197", x"1087", x"0F61", x"0DC4", x"0B68", x"07CA", x"02E1", x"FCAB",
		x"F62A", x"F07C", x"ECFE", x"EC6C", x"EEBC", x"F2B1", x"F6EC", x"FA30",
		x"FBD1", x"FBA6", x"F9F8", x"F726", x"F3CB", x"F078", x"EDA8", x"EBE2",
		x"EBB0", x"ED9A", x"F1D6", x"F808", x"FF94", x"0713", x"0D6F", x"11D5",
		x"1398", x"128F", x"0EE8", x"0932", x"024F", x"FB1D", x"F482", x"EF3B",
		x"EC88", x"ED06", x"F0F3", x"F769", x"FEE6", x"05F7", x"0BD2", x"100C",
		x"1290", x"13AC", x"13C4", x"1335", x"11FE", x"1016", x"0CFD", x"08C6",
		x"035F", x"FD66", x"F75D", x"F1FA", x"EE08", x"EC08", x"ECA2", x"F02F",
		x"F699", x"FEB6", x"073C", x"0E34", x"1256", x"1318", x"10F2", x"0D86",
		x"0AC3", x"0A21", x"0BDB", x"0F29", x"1257", x"13A8", x"11F2", x"0D2F",
		x"0636", x"FE81", x"F778", x"F1EE", x"EE63", x"EC9A", x"EBFA", x"EBC4",
		x"EC09", x"ECCD", x"EE42", x"F0F6", x"F53A", x"FB39", x"0268", x"09DA",
		x"0FDB", x"12E7", x"1232", x"0D99", x"0649", x"FDF3", x"F62E", x"F02D",
		x"EC5E", x"EA9C", x"EA65", x"EAEE", x"EB48", x"EB3D", x"EAD2", x"EAA7",
		x"EB52", x"ED57", x"F117", x"F69E", x"FDAD", x"055C", x"0C50", x"1186",
		x"141E", x"1459", x"12FC", x"1105", x"0F83", x"0F02", x"0F9E", x"10EA",
		x"125B", x"13C0", x"1476", x"13BE", x"10B7", x"0B00", x"0352", x"FB40",
		x"F401", x"EEB1", x"EB87", x"EA36", x"EA17", x"EA7C", x"EADC", x"EB96",
		x"ECCA", x"EE46", x"EF67", x"EFB7", x"EF16", x"EDA5", x"EC74", x"ECBE",
		x"EFC7", x"F5D5", x"FDE2", x"05E7", x"0C3C", x"1041", x"126F", x"1378",
		x"1411", x"1483", x"14E4", x"14F8", x"148D", x"1302", x"0F5C", x"0983",
		x"0211", x"FA31", x"F35E", x"EE7F", x"EBEB", x"EB54", x"EC65", x"EE1D",
		x"EFFC", x"F190", x"F300", x"F490", x"F665", x"F846", x"FA0D", x"FBA2",
		x"FD5A", x"FF76", x"0211", x"0540", x"08D4", x"0C87", x"0FDE", x"1293",
		x"13BF", x"12A4", x"0EC0", x"0858", x"009F", x"F8F2", x"F27A", x"EE00",
		x"EBF6", x"EC98", x"EFC7", x"F529", x"FC14", x"03A3", x"0AD9", x"104E",
		x"1361", x"13B0", x"1187", x"0D3F", x"0716", x"FF9E", x"F7D3", x"F151",
		x"ED60", x"ED17", x"F084", x"F6CF", x"FE5A", x"053A", x"097D", x"09E8",
		x"0613", x"FF18", x"F6F4", x"F092", x"ED54", x"ED07", x"EE32", x"EF15",
		x"EEE1", x"EDED", x"ED7F", x"EF27", x"F3BA", x"FAB4", x"0214", x"077A",
		x"093B", x"0720", x"01D9", x"FB07", x"F421", x"EF17", x"ED3C", x"EF63",
		x"F53D", x"FD3D", x"0585", x"0C75", x"1143", x"13B1", x"13EA", x"11EB",
		x"0E64", x"0A1D", x"05F5", x"0270", x"FF95", x"FD77", x"FBD6", x"FA77",
		x"F8BC", x"F6B3", x"F477", x"F20B", x"EFE0", x"EDD3", x"EC25", x"EB11",
		x"EAB8", x"EAA7", x"EAAC", x"EACC", x"EB00", x"EB81", x"EC86", x"EE38",
		x"F10A", x"F4EB", x"FA23", x"002B", x"0691", x"0C76", x"1121", x"1387",
		x"12C6", x"0E85", x"077C", x"FEB9", x"F620", x"EFA1", x"EC93", x"ECC3",
		x"EEA5", x"F020", x"F036", x"EEF9", x"ED99", x"ED9A", x"F01E", x"F55B",
		x"FC3E", x"02C0", x"06BD", x"0723", x"0418", x"FE80", x"F7D7", x"F1BF",
		x"EDC3", x"ED70", x"F18D", x"F95A", x"02E1", x"0B8A", x"116F", x"13F1",
		x"13C9", x"1224", x"1064", x"0FD2", x"1098", x"124C", x"1320", x"11AE",
		x"0D07", x"05F3", x"FE5A", x"F832", x"F4B8", x"F3EC", x"F566", x"F88A",
		x"FCE5", x"01A2", x"05FA", x"0985", x"0BF9", x"0DBE", x"0EF8", x"0FF2",
		x"10E3", x"11E9", x"12E1", x"13AC", x"13A7", x"1223", x"0E67", x"0860",
		x"0099", x"F8AE", x"F212", x"EDD1", x"EBBF", x"EB42", x"EBDE", x"ED05",
		x"EE55", x"EFB4", x"F0CA", x"F1A7", x"F31D", x"F552", x"F8A4", x"FCDC",
		x"0182", x"05BF", x"08EA", x"0AA1", x"0A6F", x"07DF", x"0294", x"FB41",
		x"F3C6", x"EE71", x"ECBD", x"EDFB", x"F042", x"F18F", x"F0F0", x"EF13",
		x"EDAE", x"EE95", x"F2C8", x"F964", x"0073", x"059B", x"075A", x"0530",
		x"FFF4", x"F916", x"F266", x"EDFE", x"ED1F", x"F028", x"F6B4", x"FF39",
		x"07F7", x"0ED8", x"12FF", x"13E9", x"1289", x"101A", x"0DD9", x"0C9D",
		x"0CC2", x"0E32", x"1032", x"1262", x"13F7", x"14C9", x"1523", x"1527",
		x"1507", x"14A4", x"13D2", x"1274", x"10CF", x"0EFD", x"0D99", x"0CC8",
		x"0CA5", x"0D29", x"0E12", x"0F6B", x"1114", x"12D0", x"141C", x"146F",
		x"12DA", x"0F11", x"08F3", x"0173", x"F9B6", x"F306", x"EE37", x"EBB5",
		x"EB37", x"EC49", x"EE42", x"F085", x"F298", x"F447", x"F561", x"F599",
		x"F4F8", x"F3B4", x"F231", x"F08C", x"EED2", x"ED25", x"EBE5", x"EB2B",
		x"EA9F", x"EA6E", x"EA85", x"EAD2", x"EB46", x"EC0C", x"EDAC", x"F0AE",
		x"F580", x"FC07", x"03AF", x"0B0E", x"10B9", x"1349", x"12E7", x"10A7",
		x"0E47", x"0D4F", x"0E71", x"10DE", x"1326", x"1321", x"0FED", x"09BC",
		x"0201", x"FA4F", x"F40A", x"EFBE", x"ED5A", x"EC69", x"EC0C", x"EBBF",
		x"EB66", x"EB26", x"EB3B", x"EB7D", x"EBD2", x"EC1B", x"ECB9", x"EE09",
		x"F0AF", x"F4EF", x"FAA2", x"0160", x"0878", x"0EAD", x"1293", x"13A2",
		x"11DC", x"0EA8", x"0B7D", x"09D4", x"0A26", x"0C1A", x"0EBC", x"1121",
		x"12FE", x"147D", x"1528", x"1434", x"10EC", x"0AF5", x"0334", x"FB0C",
		x"F360", x"EDB4", x"EA84", x"E99D", x"EA2B", x"EB12", x"EC19", x"ED2A",
		x"EEB3", x"F07B", x"F160", x"F0E0", x"EF47", x"EDAB", x"ED6C", x"EFBA",
		x"F4C6", x"FBBB", x"0304", x"08CC", x"0C20", x"0D3E", x"0C62", x"0A22",
		x"06D5", x"02E2", x"FEFE", x"FB57", x"F82E", x"F558", x"F311", x"F106",
		x"EF68", x"EE0F", x"ECF4", x"EC19", x"EB90", x"EB44", x"EB2A", x"EB83",
		x"EC13", x"ECDE", x"EDEC", x"EF30", x"F0B9", x"F24C", x"F447", x"F69B",
		x"F952", x"FC39", x"FF58", x"023B", x"04FE", x"0753", x"092F", x"0AAE",
		x"0BF5", x"0D31", x"0E8D", x"103D", x"1244", x"13B1", x"1397", x"10CD",
		x"0B0B", x"034C", x"FB2E", x"F427", x"EF1F", x"EC6F", x"EC1A", x"EE03",
		x"F20B", x"F83F", x"0025", x"089A", x"0FA7", x"135E", x"1320", x"0F64",
		x"0958", x"023B", x"FB13", x"F4A8", x"EF8B", x"EC7D", x"EC08", x"EE4E",
		x"F30F", x"F98D", x"00FE", x"0856", x"0E77", x"1273", x"13CC", x"1206",
		x"0D0E", x"05A3", x"FD23", x"F53D", x"EF7B", x"EC24", x"EACF", x"EA84",
		x"EAA8", x"EAD8", x"EB25", x"EC04", x"ED4F", x"EEAD", x"EF97", x"EF6E",
		x"EE5C", x"ECF2", x"EC77", x"EE1B", x"F2AC", x"F9F7", x"0273", x"0A80",
		x"1065", x"1388", x"13D6", x"1173", x"0CC7", x"0641", x"FEB7", x"F71D",
		x"F0D9", x"ECC8", x"EBF4", x"EE33", x"F2BC", x"F926", x"0030", x"06D9",
		x"0C5D", x"1060", x"12F4", x"145C", x"1505", x"1529", x"1520", x"1520",
		x"14EF", x"14C3", x"14B6", x"14B5", x"14AF", x"14BD", x"1482", x"13BF",
		x"119C", x"0D2F", x"0673", x"FE30", x"F600", x"EFAE", x"EC3C", x"EB7A",
		x"EC29", x"ECF2", x"ECD6", x"EC2A", x"EBC0", x"ED37", x"F168", x"F888",
		x"016B", x"0A02", x"1064", x"12FD", x"11A1", x"0D04", x"0675", x"FF8A",
		x"F981", x"F4EB", x"F259", x"F1A2", x"F2BE", x"F55B", x"F8FF", x"FCF9",
		x"006D", x"0251", x"01CE", x"FE9A", x"F921", x"F2F5", x"EE59", x"ED1A",
		x"EF85", x"F413", x"F86D", x"FAEA", x"FB02", x"F8BF", x"F534", x"F187",
		x"EEA6", x"ED02", x"EC6C", x"ED59", x"F03A", x"F571", x"FC69", x"040F",
		x"0B11", x"1071", x"1379", x"13E2", x"1259", x"0F7E", x"0C64", x"0995",
		x"0770", x"0610", x"055C", x"052D", x"0579", x"0677", x"080E", x"0A35",
		x"0C52", x"0E63", x"1049", x"11F0", x"1353", x"1472", x"1525", x"155A",
		x"14F9", x"1405", x"12EE", x"11E8", x"10D8", x"0F92", x"0E18", x"0C90",
		x"0AD4", x"08C8", x"0649", x"02E2", x"FE6F", x"F90D", x"F380", x"EF00",
		x"EC7C", x"ECA1", x"EF6A", x"F46D", x"FABA", x"0148", x"0735", x"0C03",
		x"0F57", x"1158", x"1275", x"12FC", x"12EA", x"1217", x"0FD3", x"0BF1",
		x"0631", x"FF09", x"F771", x"F0CB", x"ECD8", x"EC67", x"EF66", x"F4D0",
		x"FB97", x"0295", x"0919", x"0E6E", x"1226", x"1348", x"1130", x"0BB1",
		x"039C", x"FAD1", x"F324", x"EDFD", x"EB62", x"EA64", x"EA59", x"EA94",
		x"EB7C", x"EDB1", x"F22A", x"F920", x"01B8", x"09E2", x"0FFC", x"1364",
		x"14DD", x"1549", x"153B", x"14E0", x"145F", x"13BE", x"1271", x"0FA1",
		x"0A62", x"02B5", x"F9F1", x"F241", x"ED67", x"EB63", x"EB77", x"EBDD",
		x"EBD2", x"EBC3", x"ECFA", x"F075", x"F6B2", x"FF02", x"077A", x"0E5B",
		x"127C", x"144B", x"14C4", x"14A5", x"14BF", x"14D6", x"14CC", x"13F3",
		x"116C", x"0C57", x"04AF", x"FBE4", x"F400", x"EE7F", x"EB8F", x"EA78",
		x"EA3B", x"EA57", x"EADF", x"ECC1", x"F0C7", x"F74D", x"FFA9", x"0816",
		x"0EFB", x"1348", x"153F", x"156C", x"146E", x"1307", x"11CD", x"117E",
		x"122D", x"1351", x"13C1", x"126A", x"0E4E", x"07CC", x"FFEE", x"F86B",
		x"F298", x"EFA2", x"F00A", x"F3A9", x"F9EB", x"0183", x"093F", x"0F62",
		x"1309", x"13A1", x"1169", x"0D66", x"08BF", x"04A8", x"0183", x"FFC5",
		x"FF69", x"008D", x"036F", x"07DF", x"0CEB", x"1109", x"12ED", x"11A0",
		x"0D9B", x"0864", x"03AD", x"009A", x"FFB6", x"00CA", x"0331", x"0688",
		x"0A0A", x"0D81", x"1061", x"1286", x"13F0", x"14A1", x"149D", x"142C",
		x"1398", x"1343", x"1375", x"1422", x"1476", x"136A", x"1009", x"0A39",
		x"02B0", x"FA93", x"F3C5", x"EF25", x"ED00", x"ECBB", x"EDAD", x"EFBD",
		x"F2D5", x"F6D5", x"FAF3", x"FE76", x"017C", x"03E2", x"05DA", x"0767",
		x"089B", x"0A0E", x"0C46", x"0F37", x"1205", x"136B", x"1259", x"0E70",
		x"0825", x"0095", x"F95D", x"F3A6", x"F03E", x"EED6", x"EF2E", x"F0C5",
		x"F34F", x"F639", x"F977", x"FC66", x"FE98", x"FFBF", x"FFEC", x"FF48",
		x"FDBA", x"FB67", x"F83D", x"F497", x"F0D0", x"EDB8", x"EC56", x"ED94",
		x"F1D7", x"F86D", x"001E", x"0732", x"0C75", x"0EFB", x"0DD3", x"093D",
		x"0207", x"F9E8", x"F2CD", x"EE12", x"EC12", x"EC44", x"ED94", x"EEB4",
		x"EEA1", x"ED88", x"EC0D", x"EB23", x"EB13", x"EBE0", x"ED6E", x"EF9C",
		x"F258", x"F56B", x"F889", x"FAFF", x"FCA7", x"FCD3", x"FB33", x"F7E6",
		x"F365", x"EF1E", x"ECFD", x"EE2E", x"F260", x"F82B", x"FD8B", x"011B",
		x"0245", x"00E4", x"FD7D", x"F91E", x"F4E2", x"F1B0", x"EFC8", x"EF22",
		x"F004", x"F246", x"F5AB", x"F9EA", x"FE0D", x"010D", x"020D", x"0070",
		x"FC7B", x"F6E9", x"F150", x"ED78", x"ECBD", x"EF39", x"F39F", x"F818",
		x"FB0E", x"FBE4", x"FA7B", x"F7B6", x"F44A", x"F11A", x"EEBF", x"ED5E",
		x"ECB6", x"ECD3", x"ED8E", x"EED8", x"F0B1", x"F319", x"F5F3", x"F8FB",
		x"FBFA", x"FF12", x"0250", x"05AE", x"08E8", x"0B8E", x"0DAB", x"0F19",
		x"0FE0", x"0FAC", x"0E87", x"0C65", x"0972", x"062D", x"0305", x"0043",
		x"FE3B", x"FD62", x"FDAB", x"FF40", x"01A0", x"0457", x"0720", x"09FB",
		x"0CB1", x"0F21", x"1130", x"12BF", x"13EB", x"1469", x"1471", x"1432",
		x"1432", x"147A", x"14AC", x"13DF", x"1161", x"0CDB", x"0651", x"FEA7",
		x"F707", x"F0EF", x"ECE9", x"EB0F", x"EA6F", x"EAC4", x"EB93", x"EC9E",
		x"ED9D", x"EE85", x"EF6B", x"F0AF", x"F21E", x"F3BD", x"F572", x"F7BD",
		x"FABC", x"FE8B", x"0320", x"083B", x"0D61", x"119A", x"13B0", x"12F4",
		x"0F51", x"09AF", x"031B", x"FC9F", x"F6DF", x"F231", x"EED9", x"ECD8",
		x"EBDD", x"EBA9", x"EBF2", x"ECDB", x"EEEA", x"F27D", x"F7C6", x"FE68",
		x"05B0", x"0C6B", x"114D", x"12F4", x"109B", x"0A7A", x"01F7", x"F8F9",
		x"F1AF", x"ED11", x"EADF", x"EA2F", x"EA53", x"EB65", x"EE20", x"F2F8",
		x"F9D0", x"01E1", x"09E9", x"101D", x"1362", x"1346", x"1037", x"0A81",
		x"02DC", x"FA67", x"F2B0", x"ED67", x"EB17", x"EB7E", x"ED75", x"EF76",
		x"F0BF", x"F16B", x"F241", x"F41E", x"F7A1", x"FCD2", x"0336", x"09E4",
		x"0F90", x"12DC", x"1310", x"10BE", x"0D1E", x"09C2", x"0766", x"06D0",
		x"07C3", x"0A0D", x"0D18", x"100E", x"1255", x"13D3", x"1499", x"14C7",
		x"14B7", x"14B3", x"1495", x"1429", x"1306", x"10C6", x"0CAF", x"064C",
		x"FE21", x"F5E3", x"EF90", x"EC7D", x"EC19", x"ED37", x"EDF7", x"EDC5",
		x"ECDB", x"EC7C", x"EE2D", x"F2F1", x"FA65", x"02E7", x"0A75", x"0FC2",
		x"12A2", x"13D0", x"141C", x"1431", x"148E", x"14FE", x"14FB", x"13A5",
		x"0FEB", x"0977", x"0121", x"F8B3", x"F1D8", x"ED22", x"EA6F", x"E967",
		x"E9F6", x"EC86", x"F0FD", x"F762", x"FF4D", x"07AA", x"0ED5", x"1397",
		x"1563", x"151A", x"13A0", x"1164", x"0E63", x"0B16", x"0890", x"07E2",
		x"096D", x"0C84", x"0FEA", x"11D2", x"10BF", x"0C77", x"063E", x"0057",
		x"FD23", x"FDCD", x"0206", x"0838", x"0E46", x"1241", x"1303", x"10A5",
		x"0BFD", x"064A", x"00AC", x"FC18", x"F87D", x"F5DD", x"F423", x"F345",
		x"F322", x"F3C3", x"F511", x"F714", x"F9A5", x"FC8B", x"FF7C", x"020F",
		x"03FB", x"052B", x"0563", x"046C", x"028D", x"000F", x"FD2C", x"FA1D",
		x"F719", x"F45B", x"F1AB", x"EF4F", x"ED4A", x"EBC3", x"EAE8", x"EAA4",
		x"EA82", x"EA72", x"EABA", x"EC1F", x"EF7C", x"F52F", x"FCA3", x"04DD",
		x"0C2C", x"116F", x"144F", x"153F", x"1503", x"1430", x"12D5", x"10C1",
		x"0E57", x"0BF0", x"09FA", x"08D2", x"08B4", x"0975", x"0AE3", x"0CE9",
		x"0F66", x"11DC", x"139E", x"1416", x"1295", x"0F01", x"09A4", x"02D7",
		x"FB73", x"F499", x"EF59", x"EC45", x"EB44", x"EBD9", x"ED2F", x"EECD",
		x"F048", x"F170", x"F220", x"F22B", x"F1AB", x"F0C7", x"EFA9", x"EE79",
		x"ED62", x"EC4E", x"EB67", x"EAFE", x"EB25", x"EBF5", x"ED88", x"EFE6",
		x"F2C7", x"F59B", x"F765", x"F751", x"F568", x"F24C", x"EF3D", x"ED83",
		x"EE6D", x"F2A2", x"F8EF", x"FF9B", x"0423", x"0505", x"01E6", x"FC1E",
		x"F560", x"EFDC", x"ECF5", x"ED67", x"F0BD", x"F61B", x"FC25", x"01C2",
		x"0630", x"093E", x"0B3C", x"0C26", x"0BB4", x"0983", x"0542", x"FF70",
		x"F906", x"F2FD", x"EEA5", x"ECB3", x"ED79", x"F09E", x"F505", x"F9F2",
		x"FE64", x"020C", x"04D5", x"06C8", x"07E9", x"0816", x"0775", x"05AC",
		x"0312", x"FFBD", x"FC31", x"F8FB", x"F696", x"F5A1", x"F696", x"FA09",
		x"FFA1", x"068F", x"0D18", x"1183", x"131C", x"11CF", x"0F01", x"0C29",
		x"0A72", x"0A5A", x"0B95", x"0DB6", x"1060", x"12ED", x"14A8", x"14C3",
		x"12AA", x"0E16", x"07AF", x"0004", x"F87C", x"F21C", x"EDA0", x"EB82",
		x"EB6C", x"ECBE", x"EEAF", x"F095", x"F225", x"F35A", x"F3EF", x"F3CD",
		x"F2F9", x"F1DB", x"F07F", x"EF0B", x"ED7C", x"EC0D", x"EB2D", x"EABE",
		x"EAB6", x"EABA", x"EAC7", x"EAF7", x"EBA0", x"ECED", x"EF17", x"F25C",
		x"F6BC", x"FC0A", x"0224", x"085E", x"0DEB", x"1208", x"13DC", x"127C",
		x"0DBB", x"065C", x"FDFC", x"F62F", x"F025", x"EC77", x"EB3D", x"EC60",
		x"EF6C", x"F3A3", x"F870", x"FD11", x"010B", x"03FF", x"0619", x"0756",
		x"07C5", x"07CD", x"0757", x"06C0", x"05EF", x"04C2", x"02C6", x"FFE0",
		x"FBE9", x"F70C", x"F236", x"EEA1", x"ED7A", x"EFA4", x"F4B7", x"FB7C",
		x"021D", x"06DF", x"0801", x"0502", x"FEA9", x"F6F9", x"F099", x"ED53",
		x"ED2B", x"EEB9", x"F042", x"F05A", x"EF08", x"ED9B", x"EE23", x"F219",
		x"F90D", x"00F4", x"0767", x"0AE3", x"0B23", x"08D6", x"04FF", x"0061",
		x"FBE1", x"F890", x"F767", x"F933", x"FDDC", x"049F", x"0B97", x"10F9",
		x"1318", x"123D", x"0F8A", x"0C68", x"0A7A", x"0A4E", x"0BFD", x"0EB0",
		x"1174", x"136E", x"1486", x"14D3", x"14C9", x"14A4", x"145C", x"13BE",
		x"128B", x"109B", x"0DF7", x"0B0C", x"081C", x"0527", x"0205", x"FEDB",
		x"FBE8", x"F946", x"F747", x"F5D6", x"F503", x"F518", x"F600", x"F79B",
		x"F9CC", x"FC9E", x"000B", x"03BB", x"0742", x"0A37", x"0CB2", x"0EAA",
		x"1049", x"1177", x"1271", x"1344", x"1415", x"14C0", x"14DE", x"1431",
		x"12D1", x"10D7", x"0EDB", x"0DB0", x"0DB3", x"0EF3", x"10E6", x"12CA",
		x"1377", x"11C4", x"0D2A", x"0657", x"FEAD", x"F7E0", x"F2BF", x"EF8A",
		x"ED93", x"EC7C", x"EBD2", x"EB2C", x"EABF", x"EAA8", x"EB7A", x"EDC4",
		x"F209", x"F828", x"FF70", x"0720", x"0DDB", x"126A", x"13D4", x"11DE",
		x"0CF0", x"062C", x"FEB2", x"F794", x"F1C6", x"EDF2", x"EC21", x"EBF2",
		x"ED2D", x"EF68", x"F217", x"F495", x"F67D", x"F730", x"F68D", x"F47C",
		x"F1B8", x"EEAB", x"ECB0", x"ECBD", x"EF81", x"F510", x"FCBC", x"050C",
		x"0C8C", x"121C", x"14B7", x"1483", x"11C5", x"0CFD", x"064E", x"FE7D",
		x"F691", x"F059", x"ED71", x"EE83", x"F2D4", x"F8C4", x"FE62", x"01EB",
		x"023E", x"FF38", x"F9B9", x"F39E", x"EEFF", x"ED17", x"EDFF", x"F0C3",
		x"F45E", x"F78F", x"F99E", x"F9E5", x"F874", x"F59A", x"F224", x"EECC",
		x"EC76", x"EC2A", x"EEA1", x"F40A", x"FB5D", x"0323", x"09FF", x"0F2F",
		x"1272", x"1394", x"127E", x"0EFD", x"0913", x"015C", x"F913", x"F1B6",
		x"ECE6", x"EB62", x"EC8B", x"EED5", x"F0D8", x"F219", x"F2B6", x"F367",
		x"F4AF", x"F6D2", x"F9F7", x"FDF0", x"027F", x"06FB", x"0AB8", x"0D35",
		x"0E49", x"0DBD", x"0B6C", x"0720", x"010B", x"F9ED", x"F324", x"EE55",
		x"EC4B", x"ECD7", x"EFA7", x"F3D9", x"F8D2", x"FDCD", x"0205", x"0517",
		x"068B", x"0658", x"0435", x"001A", x"FA4C", x"F414", x"EEFF", x"ECCF",
		x"EDE2", x"F116", x"F468", x"F5B5", x"F443", x"F0F0", x"EE0D", x"ED92",
		x"F0BF", x"F6C6", x"FD6E", x"02A8", x"0502", x"046E", x"0176", x"FD32",
		x"F897", x"F4BC", x"F234", x"F1B6", x"F3BF", x"F860", x"FF1E", x"0686",
		x"0D64", x"11F0", x"13AB", x"1299", x"0F92", x"0BD1", x"0851", x"058C",
		x"0381", x"01F9", x"0080", x"FE99", x"FC17", x"F91D", x"F602", x"F2F4",
		x"F02E", x"EE02", x"EC9E", x"EBFE", x"EBE5", x"EC26", x"ECDB", x"EDEA",
		x"EF88", x"F1A2", x"F42E", x"F6BE", x"F8C2", x"F9E5", x"FA29", x"F998",
		x"F83E", x"F5E6", x"F322", x"F043", x"EDC3", x"EBF9", x"EB73", x"ECC4",
		x"F00A", x"F560", x"FC08", x"036A", x"0A94", x"104B", x"132A", x"1243",
		x"0DD3", x"06D8", x"FF00", x"F7D9", x"F254", x"EEAB", x"ECC7", x"EC50",
		x"ECCB", x"EDD7", x"EF86", x"F1BE", x"F4AF", x"F827", x"FBAC", x"FED2",
		x"014C", x"0305", x"044E", x"0597", x"0793", x"0A86", x"0E3E", x"11A7",
		x"1320", x"11B3", x"0D50", x"06AB", x"FF34", x"F8A2", x"F41C", x"F2E0",
		x"F570", x"FB63", x"030E", x"0AB5", x"107E", x"1373", x"13CB", x"1291",
		x"1142", x"10F8", x"11D0", x"131B", x"13E4", x"13F5", x"13F3", x"144B",
		x"1491", x"13BA", x"107A", x"0A85", x"02A5", x"FA47", x"F30B", x"EE48",
		x"ECFB", x"EF41", x"F4AC", x"FC31", x"0459", x"0BBA", x"111D", x"140E",
		x"14F3", x"1496", x"1449", x"1456", x"149F", x"1467", x"138C", x"1270",
		x"1177", x"1142", x"11C3", x"12CA", x"13ED", x"148E", x"14C1", x"1476",
		x"1435", x"1408", x"1438", x"1497", x"1511", x"1525", x"14EB", x"13F6",
		x"1283", x"10DA", x"0EF2", x"0CBD", x"0A03", x"06F0", x"03F0", x"0154",
		x"FF80", x"FE8F", x"FED4", x"0055", x"02E6", x"0604", x"0920", x"0C10",
		x"0E4C", x"0FEA", x"1065", x"0FB6", x"0E32", x"0BFE", x"0953", x"0636",
		x"0342", x"00CA", x"FF44", x"FEC7", x"FF27", x"0061", x"0263", x"053E",
		x"088D", x"0C10", x"0F8E", x"126D", x"13CA", x"12F5", x"0F6E", x"09C2",
		x"02D2", x"FBCC", x"F56B", x"F082", x"ED38", x"EB5B", x"EA8D", x"EA6F",
		x"EA7B", x"EAD7", x"EB8A", x"EC56", x"ED80", x"EED8", x"F087", x"F2B3",
		x"F567", x"F84F", x"FB33", x"FDF7", x"0049", x"0225", x"035C", x"0451",
		x"0593", x"07B3", x"0AD9", x"0E85", x"11EE", x"138C", x"1245", x"0DDD",
		x"0766", x"000C", x"F95F", x"F44E", x"F1BF", x"F210", x"F523", x"FA59",
		x"0124", x"0891", x"0F04", x"1285", x"11D4", x"0CE9", x"0513", x"FC2F",
		x"F435", x"EE90", x"EBB0", x"EAF2", x"EB2F", x"EB64", x"EB6E", x"EB92",
		x"ECC8", x"F028", x"F66F", x"FEEE", x"07DE", x"0F13", x"12CD", x"127F",
		x"0E7F", x"0820", x"00DB", x"FA05", x"F49C", x"F0F8", x"EF60", x"EF90",
		x"F143", x"F3E9", x"F743", x"FAD8", x"FDC5", x"FF22", x"FE44", x"FAAD",
		x"F56C", x"F064", x"ED6F", x"EDCE", x"F16F", x"F70F", x"FCFD", x"021F",
		x"05C3", x"081C", x"09C7", x"0B11", x"0C94", x"0E72", x"10C0", x"12E8",
		x"13E3", x"12C1", x"0EC0", x"0863", x"00BD", x"F94C", x"F2FB", x"EE71",
		x"EBBE", x"EAAC", x"EAAC", x"EB3F", x"EBEB", x"EC73", x"ECA5", x"EC86",
		x"EC6F", x"EC4E", x"EC1E", x"EBC3", x"EB63", x"EB3D", x"EBD6", x"ED80",
		x"F0B1", x"F58B", x"FBE7", x"0311", x"0A2E", x"1011", x"1394", x"13E1",
		x"1106", x"0B97", x"04BB", x"FD70", x"F689", x"F0DA", x"ED19", x"EC0C",
		x"EDEA", x"F27C", x"F914", x"00B0", x"082A", x"0E69", x"129E", x"1496",
		x"1461", x"125C", x"0F20", x"0B40", x"0748", x"03B5", x"0121", x"0022",
		x"010D", x"03FD", x"0890", x"0D8F", x"1153", x"120B", x"0F52", x"0A51",
		x"0591", x"0369", x"04B6", x"0906", x"0E41", x"11DC", x"1232", x"0F2D",
		x"0A85", x"06B1", x"054E", x"0715", x"0B51", x"1011", x"130A", x"1292",
		x"0E5A", x"06E0", x"FDE8", x"F52D", x"EED0", x"EBD4", x"EC42", x"EF3C",
		x"F3A8", x"F888", x"FCAD", x"FF63", x"001E", x"FF28", x"FCF3", x"F9FE",
		x"F6A4", x"F2FE", x"EFB5", x"ED24", x"EBA6", x"EAE9", x"EAA3", x"EA86",
		x"EAAE", x"EB1F", x"EB9C", x"EBEA", x"EBFF", x"EBD1", x"EB6C", x"EAF1",
		x"EAB4", x"EB34", x"ECD3", x"EFEB", x"F49F", x"FABA", x"01D2", x"08AF",
		x"0E84", x"128F", x"1458", x"13BA", x"1104", x"0CBA", x"07F7", x"0388",
		x"FFDE", x"FD81", x"FCC4", x"FE30", x"0189", x"0678", x"0BEB", x"1091",
		x"1322", x"12D0", x"0FC2", x"0B36", x"06AB", x"0333", x"018D", x"01CE",
		x"03B0", x"0696", x"0A33", x"0E0C", x"116C", x"134F", x"12BA", x"0F08",
		x"08C0", x"0122", x"F992", x"F34E", x"EF57", x"EE15", x"EFC8", x"F415",
		x"FA91", x"0250", x"0A0C", x"104C", x"13BB", x"1412", x"122C", x"0F69",
		x"0CE2", x"0AE4", x"094A", x"07B6", x"05F9", x"03D7", x"01CA", x"FFF0",
		x"FE59", x"FCB0", x"FAA1", x"F812", x"F507", x"F1DF", x"EECA", x"EC96",
		x"EC28", x"EE35", x"F2CF", x"F979", x"00E9", x"0802", x"0DCC", x"11CF",
		x"141D", x"1508", x"14E0", x"1430", x"138E", x"1397", x"1434", x"1496",
		x"135B", x"0FC8", x"09A1", x"01D1", x"F997", x"F27D", x"EDEC", x"ECE4",
		x"EFA2", x"F5C1", x"FDEF", x"0649", x"0D58", x"1237", x"14E3", x"161C",
		x"15A5", x"1388", x"0F73", x"0965", x"01E7", x"F9DD", x"F2CE", x"EE16",
		x"ECDC", x"EF2A", x"F477", x"FBB0", x"03B2", x"0B43", x"10FB", x"13D0",
		x"13C9", x"11EE", x"0F86", x"0D92", x"0C20", x"0ADA", x"0953", x"0784",
		x"0539", x"028E", x"FF93", x"FC36", x"F8F5", x"F606", x"F39E", x"F200",
		x"F111", x"F0DB", x"F18A", x"F2FF", x"F54D", x"F822", x"FB78", x"FED3",
		x"01ED", x"04E0", x"0767", x"0975", x"0B02", x"0C3A", x"0D8E", x"0F74",
		x"11E3", x"13E3", x"142A", x"1185", x"0BFF", x"0474", x"FC8C", x"F575",
		x"F041", x"ED69", x"ED61", x"F02E", x"F5B4", x"FD13", x"0530", x"0C85",
		x"11E1", x"14CC", x"155A", x"14C4", x"1435", x"1451", x"14E8", x"151D",
		x"140B", x"11AD", x"0E06", x"0912", x"0301", x"FC73", x"F607", x"F0B4",
		x"ED4E", x"ECAF", x"EF46", x"F4BF", x"FC69", x"04C6", x"0C6A", x"11BC",
		x"1429", x"141A", x"12AE", x"111A", x"107F", x"1101", x"124F", x"13B7",
		x"147A", x"14B8", x"14C1", x"14D1", x"14DB", x"14F1", x"14B4", x"1414",
		x"12ED", x"11AD", x"10E5", x"10F4", x"11DA", x"1324", x"13EF", x"1306",
		x"0F85", x"0954", x"0140", x"F8E2", x"F1D6", x"ED87", x"EC9C", x"EF32",
		x"F453", x"FB0A", x"01D2", x"079A", x"0BA0", x"0D63", x"0D0E", x"0B14",
		x"0828", x"0476", x"00C9", x"FD9D", x"FBA2", x"FB14", x"FC1C", x"FE7F",
		x"01E1", x"05C3", x"096B", x"0C62", x"0E03", x"0E2D", x"0CC2", x"0A0B",
		x"067B", x"0251", x"FE55", x"FB70", x"FA56", x"FBCA", x"FFD4", x"05D8",
		x"0C5C", x"116D", x"1392", x"127F", x"0F41", x"0B5D", x"0878", x"07A4",
		x"08CD", x"0B6C", x"0E8B", x"1176", x"137F", x"148E", x"14D1", x"145C",
		x"136D", x"11F0", x"0FFC", x"0DA8", x"0B61", x"0985", x"0888", x"088A",
		x"096F", x"0B3B", x"0D42", x"0F7B", x"1170", x"130F", x"1429", x"14CC",
		x"14F2", x"149E", x"13C5", x"1291", x"1148", x"1051", x"0FB8", x"0F6C",
		x"0F88", x"1033", x"1159", x"12CA", x"13F8", x"14A9", x"14E1", x"14C7",
		x"1421", x"12FB", x"115F", x"0F8A", x"0D9A", x"0BCB", x"0A45", x"094E",
		x"08F0", x"0929", x"09E9", x"0B25", x"0CE7", x"0F05", x"112F", x"1321",
		x"140A", x"1328", x"0FD8", x"0A17", x"02BB", x"FAEA", x"F3D3", x"EE95",
		x"EBB3", x"EACA", x"EB06", x"EBA7", x"EC48", x"ECEF", x"EDED", x"EF8E",
		x"F208", x"F5F8", x"FBC2", x"0309", x"0A78", x"1050", x"1368", x"133F",
		x"10B4", x"0D10", x"096A", x"06B2", x"0511", x"0401", x"02C8", x"00B2",
		x"FD26", x"F849", x"F2ED", x"EEB2", x"ED03", x"EE84", x"F2DE", x"F8F4",
		x"FEF0", x"02BC", x"032D", x"0038", x"FB1F", x"F548", x"F043", x"ED8E",
		x"EE35", x"F26C", x"F960", x"018B", x"0953", x"0F4F", x"1312", x"145A",
		x"1313", x"0F82", x"09DB", x"02A6", x"FB19", x"F43B", x"EF12", x"EC36",
		x"EC19", x"EEC9", x"F3FD", x"FB08", x"02DE", x"0A35", x"1011", x"1393",
		x"143F", x"124E", x"0E73", x"0992", x"0467", x"FF7A", x"FB3C", x"F7E6",
		x"F5C6", x"F4BB", x"F4CB", x"F641", x"F9A0", x"FEC5", x"051E", x"0B6A",
		x"1063", x"12BD", x"120B", x"0E24", x"07EF", x"0096", x"F92E", x"F2D2",
		x"EE6B", x"EC83", x"ED24", x"F045", x"F56C", x"FC07", x"0351", x"0A61",
		x"101F", x"1398", x"1442", x"11D2", x"0CA4", x"057B", x"FD4A", x"F594",
		x"EF8B", x"EC45", x"EBAF", x"ED27", x"EF8D", x"F1C9", x"F330", x"F3A3",
		x"F2F9", x"F15F", x"EF3C", x"ED08", x"EBB0", x"EC12", x"EF18", x"F4E9",
		x"FCAA", x"04E1", x"0BE6", x"10EC", x"13BC", x"1501", x"14D5", x"1365",
		x"102C", x"0A85", x"02A4", x"F9D1", x"F231", x"EDA8", x"ED36", x"F076",
		x"F626", x"FD18", x"0420", x"0A58", x"0F5A", x"1295", x"13FB", x"13AE",
		x"121C", x"0FD3", x"0D80", x"0BB4", x"0AE6", x"0B77", x"0D40", x"0FE4",
		x"1260", x"13AF", x"12C9", x"0F59", x"098F", x"0275", x"FB1E", x"F4D7",
		x"F039", x"ED6F", x"EBF1", x"EB41", x"EAEC", x"EAE2", x"EB0B", x"EBA4",
		x"ED09", x"EFE5", x"F480", x"FB19", x"02E6", x"0AA2", x"10A2", x"1352",
		x"1221", x"0D84", x"066D", x"FE5C", x"F6F0", x"F130", x"ED86", x"EB9B",
		x"EAF9", x"EB0B", x"EB3C", x"EB66", x"EBC2", x"ECBB", x"EEE9", x"F2A5",
		x"F7E6", x"FE55", x"054B", x"0BF6", x"10F5", x"1394", x"1352", x"10CF",
		x"0CF3", x"08E4", x"0561", x"0295", x"00C1", x"FF63", x"FDC1", x"FB4D",
		x"F7BE", x"F383", x"EF88", x"ED31", x"EDA3", x"F170", x"F79D", x"FEAB",
		x"04AC", x"082F", x"08FA", x"0752", x"040E", x"FFE6", x"FBE8", x"F88C",
		x"F68C", x"F6AF", x"F934", x"FE06", x"045D", x"0B42", x"10C7", x"137D",
		x"1281", x"0E06", x"0736", x"FF66", x"F81D", x"F22B", x"EE02", x"EBFE",
		x"EC86", x"EFC4", x"F593", x"FD22", x"0520", x"0C45", x"115D", x"13BD",
		x"1370", x"10F5", x"0D64", x"0996", x"0625", x"0345", x"00AC", x"FE2C",
		x"FB95", x"F92C", x"F74E", x"F5D4", x"F483", x"F30A", x"F19B", x"F04C",
		x"EEFC", x"ED89", x"EC33", x"EBF0", x"EDE7", x"F2C4", x"FA11", x"022B",
		x"0994", x"0F34", x"12B8", x"1442", x"13F0", x"11C4", x"0DBF", x"07D5",
		x"005A", x"F85A", x"F181", x"ED97", x"EDE0", x"F275", x"FA3A", x"032A",
		x"0B1B", x"10AA", x"13D4", x"1538", x"1567", x"13FC", x"105C", x"0A46",
		x"0292", x"FA4A", x"F2E4", x"ED57", x"EA91", x"EB01", x"EE75", x"F469",
		x"FC46", x"04B7", x"0C90", x"123E", x"153C", x"15E7", x"156A", x"1497",
		x"139D", x"123D", x"105D", x"0ECE", x"0E58", x"0F47", x"1120", x"12F7",
		x"132D", x"10BB", x"0B62", x"03F2", x"FC45", x"F5DD", x"F15D", x"EEAF",
		x"ED09", x"EC10", x"EB5E", x"EAF6", x"EAC2", x"EAE8", x"EB54", x"EC04",
		x"ED12", x"EE3A", x"EF93", x"F12E", x"F340", x"F5C8", x"F8AA", x"FBB5",
		x"FEAE", x"0192", x"043C", x"06AF", x"08DC", x"0AAF", x"0BD7", x"0C66",
		x"0C36", x"0B28", x"0913", x"0609", x"0240", x"FDFC", x"F972", x"F4C2",
		x"F07F", x"ED40", x"EBD6", x"ECB9", x"F064", x"F6B5", x"FEE3", x"0798",
		x"0EDF", x"12F3", x"1306", x"0F7E", x"09EC", x"0441", x"FFE7", x"FDD6",
		x"FEE2", x"02EF", x"08D6", x"0E79", x"1201", x"1251", x"0F6B", x"0A60",
		x"04BE", x"FFEB", x"FCA9", x"FB16", x"FA6F", x"F9CA", x"F84B", x"F559",
		x"F1A4", x"EE82", x"ED89", x"EFD3", x"F516", x"FC4D", x"03AD", x"092A",
		x"0B51", x"096A", x"0406", x"FCA1", x"F536", x"EF9D", x"EC9D", x"EC43",
		x"EDD0", x"F01A", x"F1F8", x"F28A", x"F1B4", x"EFF3", x"EDE8", x"EC37",
		x"EB90", x"ED00", x"F11C", x"F7ED", x"0037", x"0866", x"0F04", x"134A",
		x"157D", x"1636", x"15C6", x"1423", x"10E4", x"0B8C", x"0404", x"FB56",
		x"F367", x"EDCC", x"EB61", x"EB46", x"EC35", x"ED7B", x"EEA8", x"EFB5",
		x"F080", x"F0CE", x"F04F", x"EF53", x"EDD6", x"EC6A", x"EB8A", x"EB38",
		x"EB19", x"EADC", x"EAA7", x"EB00", x"ECDD", x"F08B", x"F637", x"FD8E",
		x"0577", x"0C70", x"117C", x"143E", x"14DA", x"1400", x"126C", x"10A4",
		x"0F48", x"0EC7", x"0F65", x"10E1", x"1290", x"1353", x"1209", x"0E0C",
		x"0794", x"FFE9", x"F8BD", x"F3AB", x"F140", x"F148", x"F342", x"F6AF",
		x"FAE6", x"FF24", x"0297", x"049A", x"04B9", x"030B", x"FFBA", x"FB95",
		x"F785", x"F455", x"F288", x"F22D", x"F3C2", x"F78D", x"FD9C", x"04F9",
		x"0C3B", x"1172", x"13E2", x"1341", x"1096", x"0CED", x"0951", x"0654",
		x"03FC", x"023A", x"0078", x"FE8D", x"FC6D", x"FA31", x"F7C2", x"F525",
		x"F2AD", x"F08D", x"EF06", x"EDD6", x"ECAF", x"EB98", x"EADB", x"EA9F",
		x"EB1A", x"EC47", x"EDC0", x"EF28", x"EFF0", x"EFDB", x"EF24", x"EDF4",
		x"ECA3", x"EB9E", x"EB14", x"EAD7", x"EAF6", x"EB18", x"EB63", x"EC13",
		x"EDDF", x"F159", x"F71D", x"FEBA", x"06F6", x"0E45", x"128A", x"12FB",
		x"0F68", x"089E", x"0070", x"F8BE", x"F2D1", x"EF37", x"EDDC", x"EECA",
		x"F1F1", x"F74A", x"FE43", x"0601", x"0D23", x"122F", x"145B", x"13AA",
		x"1146", x"0E9B", x"0C95", x"0B50", x"0A56", x"0921", x"0732", x"0486",
		x"0105", x"FCD5", x"F86F", x"F469", x"F17F", x"EFDB", x"EFC3", x"F168",
		x"F524", x"FB33", x"02B4", x"0A60", x"107D", x"1419", x"14FF", x"13D5",
		x"11E4", x"1047", x"0FAD", x"1044", x"1191", x"131C", x"1422", x"13FA",
		x"11E5", x"0D0F", x"0598", x"FCDB", x"F4DF", x"EEFC", x"EBAB", x"EA82",
		x"EA5F", x"EAC3", x"EC33", x"EF47", x"F4A7", x"FC19", x"0482", x"0C0D",
		x"1149", x"13C6", x"1424", x"132C", x"1159", x"0EC2", x"0B8C", x"082A",
		x"054B", x"039E", x"0345", x"041F", x"05EF", x"084F", x"0B1B", x"0E25",
		x"110D", x"134A", x"141B", x"132C", x"100B", x"0AAB", x"0390", x"FBD5",
		x"F4D7", x"EF8F", x"EC5D", x"EAFC", x"EAF9", x"EB95", x"EC59", x"ED14",
		x"ED9A", x"EDE4", x"EDE9", x"ED71", x"ECB6", x"EBCA", x"EB27", x"EAEA",
		x"EB34", x"EBB8", x"EC20", x"EC27", x"EBDB", x"EB91", x"EBCD", x"ECB5",
		x"EDCA", x"EE4F", x"EDD1", x"ECB6", x"EC7A", x"EE3C", x"F2BA", x"F93E",
		x"00EB", x"080E", x"0CF2", x"0EB3", x"0CD8", x"07FB", x"00EE", x"F942",
		x"F24F", x"EDA2", x"EC30", x"EDD3", x"F13F", x"F537", x"F8A0", x"FB5D",
		x"FD60", x"FED9", x"FFA8", x"FFDB", x"FF7D", x"FE86", x"FCFE", x"FAD6",
		x"F85E", x"F5BC", x"F311", x"F0A9", x"EE95", x"ECE0", x"EB9F", x"EB00",
		x"EAF9", x"EB57", x"EBFA", x"EC60", x"EC85", x"EC1B", x"EB49", x"EAA7",
		x"EAE0", x"EBDB", x"ECFC", x"ED92", x"ED3A", x"EC83", x"EC51", x"EDC1",
		x"F1AD", x"F814", x"000E", x"07D3", x"0DDB", x"1121", x"11B7", x"102A",
		x"0D4F", x"099D", x"05EA", x"02DF", x"013D", x"01AF", x"0475", x"0925",
		x"0E3E", x"120F", x"1313", x"10DD", x"0C03", x"05EE", x"FFE4", x"FAD6",
		x"F72F", x"F4EC", x"F35A", x"F220", x"F0D0", x"EF50", x"EDD7", x"EC82",
		x"EB8A", x"EB1C", x"EB20", x"EB77", x"EC14", x"ECBC", x"ECFF", x"ECEB",
		x"EC64", x"EBC0", x"EB45", x"EB36", x"EB98", x"EC5B", x"ED77", x"EE8D",
		x"EFC5", x"F112", x"F2B6", x"F493", x"F6D5", x"F9E0", x"FDD6", x"02B6",
		x"0827", x"0D6B", x"119E", x"13F9", x"1390", x"1028", x"0A1C", x"024D",
		x"FA00", x"F2D8", x"EE0F", x"EC67", x"EDB3", x"F12A", x"F57B", x"F97D",
		x"FCB4", x"FE9C", x"FEF0", x"FDAA", x"FB10", x"F76F", x"F354", x"EFBC",
		x"ED2E", x"EC30", x"ED1A", x"EFF6", x"F4CE", x"FB28", x"027B", x"09A3",
		x"0F6B", x"126C", x"11A9", x"0D2C", x"05F2", x"FDBE", x"F668", x"F120",
		x"EEC9", x"EFA1", x"F39F", x"FA28", x"01E3", x"0989", x"0FA5", x"136C",
		x"14B4", x"1455", x"13BC", x"13AC", x"141B", x"147F", x"1448", x"1396",
		x"130C", x"1336", x"13FD", x"14A8", x"1410", x"1100", x"0B30", x"0322",
		x"FA51", x"F2AB", x"ED9E", x"EC67", x"EEB3", x"F3F2", x"FAC2", x"01D6",
		x"082A", x"0CD7", x"0FD4", x"10FF", x"10E5", x"0F92", x"0D69", x"0A8B",
		x"071D", x"036A", x"FF76", x"FBBC", x"F834", x"F52D", x"F288", x"F0A1",
		x"EF46", x"EE52", x"EDB6", x"ED7A", x"EDC8", x"EE61", x"EF68", x"F106",
		x"F36E", x"F6D5", x"FB32", x"00D2", x"0728", x"0D6F", x"1204", x"13A8",
		x"11E1", x"0DBE", x"0921", x"05A0", x"043D", x"050C", x"07A2", x"0B05",
		x"0E77", x"1119", x"12C0", x"12D9", x"112E", x"0D12", x"068A", x"FE92",
		x"F6B4", x"F058", x"EC74", x"EB0E", x"EB4E", x"EC39", x"ECF0", x"ECB7",
		x"EBBD", x"EAE2", x"EAFA", x"EC7C", x"EFF0", x"F537", x"FC20", x"03E8",
		x"0B4E", x"10CF", x"13D8", x"146B", x"1388", x"1255", x"1199", x"11E3",
		x"12DF", x"1401", x"14C1", x"14CC", x"1425", x"1309", x"1187", x"0FD1",
		x"0E03", x"0C3C", x"0A64", x"0840", x"0603", x"0402", x"0211", x"0008",
		x"FDB6", x"FB2A", x"F879", x"F5ED", x"F348", x"F0AA", x"EE0C", x"EC47",
		x"EC72", x"EF75", x"F55B", x"FD08", x"04E6", x"0B97", x"1035", x"1300",
		x"1478", x"1538", x"1590", x"1590", x"1556", x"14A3", x"12EB", x"0F43",
		x"0942", x"0123", x"F881", x"F16E", x"ED09", x"EB3A", x"EAE9", x"EB2B",
		x"EBBC", x"ED13", x"EFF6", x"F551", x"FCCC", x"0554", x"0D07", x"11E7",
		x"127F", x"0F16", x"087B", x"00B0", x"F92D", x"F365", x"EFBE", x"EE51",
		x"EEF1", x"F190", x"F624", x"FCA1", x"044E", x"0BA8", x"10DC", x"127F",
		x"101D", x"0A8D", x"0334", x"FB80", x"F4D7", x"EFF4", x"ECF6", x"EBAA",
		x"EBEF", x"EDAF", x"F0B5", x"F47E", x"F840", x"FB09", x"FC3B", x"FB90",
		x"F917", x"F55A", x"F138", x"EDD8", x"EC74", x"EE02", x"F26B", x"F891",
		x"FF27", x"04ED", x"0980", x"0C96", x"0E6D", x"0F84", x"106B", x"119F",
		x"130A", x"142D", x"1453", x"12AA", x"0EFF", x"093B", x"01DA", x"FA0A",
		x"F319", x"EE51", x"ECE9", x"EF0C", x"F435", x"FB4B", x"02CF", x"0998",
		x"0EBB", x"120A", x"13BD", x"1477", x"1488", x"13EB", x"125E", x"0FA6",
		x"0BB2", x"06FB", x"017B", x"FB79", x"F5A7", x"F08A", x"ED2C", x"EC28",
		x"EDF5", x"F298", x"F982", x"0182", x"091D", x"0F3A", x"130C", x"1475",
		x"136A", x"0FCB", x"09D9", x"024A", x"FA40", x"F2F3", x"EE10", x"EC91",
		x"EE74", x"F253", x"F631", x"F85A", x"F88C", x"F710", x"F452", x"F13A",
		x"EE6F", x"EC89", x"EBA8", x"EBEE", x"ED75", x"F086", x"F578", x"FC25",
		x"03E1", x"0B4E", x"10DF", x"1320", x"1139", x"0B91", x"036F", x"FAE5",
		x"F3A3", x"EE89", x"EBB5", x"EA85", x"EA68", x"EB02", x"ECC1", x"F054",
		x"F64A", x"FE26", x"0671", x"0D8B", x"1248", x"1481", x"14E8", x"1444",
		x"132C", x"1203", x"1146", x"10E4", x"10AC", x"1077", x"103F", x"104C",
		x"1100", x"121E", x"1371", x"1474", x"146F", x"12D7", x"0EED", x"08EA",
		x"0168", x"F9B0", x"F2FD", x"EE2C", x"EB8F", x"EAB6", x"EB1E", x"EB96",
		x"EB9D", x"EB42", x"EB27", x"EBEE", x"EE04", x"F19A", x"F6DC", x"FDDF",
		x"0597", x"0C91", x"1161", x"1367", x"1320", x"119D", x"1014", x"0F81",
		x"1031", x"11C2", x"135B", x"1463", x"14DB", x"1512", x"1534", x"14A2",
		x"12B2", x"0E8B", x"07FB", x"FFDB", x"F7AD", x"F130", x"ED1E", x"EB6F",
		x"EB27", x"EB70", x"EBF9", x"ED07", x"EEEC", x"F200", x"F62E", x"FB9F",
		x"022E", x"0914", x"0F02", x"12DA", x"13E1", x"122F", x"0E7B", x"09AE",
		x"04A0", x"0056", x"FCF4", x"FA96", x"F8CE", x"F74E", x"F5D0", x"F44A",
		x"F29F", x"F0CD", x"EEEA", x"ED35", x"EBD3", x"EAED", x"EA7C", x"EA90",
		x"EB2D", x"EBF9", x"ECA4", x"ED5C", x"EE30", x"EFA0", x"F1FC", x"F549",
		x"F991", x"FED5", x"04B1", x"0AA0", x"0FCF", x"1319", x"1387", x"10DC",
		x"0B84", x"0458", x"FCB1", x"F59E", x"F011", x"EC8C", x"EB91", x"ED65",
		x"F225", x"F929", x"016D", x"0981", x"0FF1", x"1365", x"138D", x"1148",
		x"0E6D", x"0CDF", x"0D6C", x"0FA6", x"124A", x"13B3", x"1287", x"0DF7",
		x"0657", x"FD48", x"F4D8", x"EF1F", x"ED46", x"EF63", x"F459", x"FA87",
		x"0029", x"03AA", x"03EB", x"0095", x"FAAC", x"F403", x"EEF1", x"ECF9",
		x"EDDC", x"F03A", x"F233", x"F291", x"F108", x"EEB4", x"EDA8", x"EFBC",
		x"F567", x"FD27", x"04DF", x"0AD6", x"0E97", x"107F", x"1157", x"11DE",
		x"129A", x"137D", x"146A", x"14A8", x"1324", x"0F41", x"08E0", x"0112",
		x"F91E", x"F297", x"EE22", x"EBB6", x"EB1C", x"EB7E", x"EC6A", x"EDB9",
		x"EF4D", x"F0E4", x"F27D", x"F415", x"F577", x"F6D0", x"F810", x"F985",
		x"FB29", x"FD97", x"0130", x"05CD", x"0AB8", x"0F28", x"11FC", x"123E",
		x"0F97", x"0A71", x"03F1", x"FE23", x"FAE8", x"FB26", x"FEB4", x"045D",
		x"0ABF", x"0FFF", x"1286", x"1154", x"0CA5", x"0545", x"FD28", x"F5CE",
		x"F015", x"EC7A", x"EB10", x"EC4A", x"F063", x"F750", x"FFD6", x"0878",
		x"0F3E", x"12FC", x"1352", x"1178", x"0F45", x"0E4C", x"0F43", x"1145",
		x"12E1", x"1237", x"0E57", x"07DA", x"00AD", x"FAB8", x"F754", x"F693",
		x"F84F", x"FBD8", x"0069", x"04E1", x"080E", x"0983", x"0874", x"050A",
		x"FF65", x"F8C3", x"F286", x"EE52", x"ED2B", x"EF67", x"F4C7", x"FC4E",
		x"0488", x"0BDC", x"1126", x"13CE", x"13F2", x"11CE", x"0E27", x"09DE",
		x"05B0", x"023C", x"FF86", x"FD71", x"FB8F", x"F9AE", x"F788", x"F51D",
		x"F2B1", x"F09E", x"EEDA", x"ED60", x"EC27", x"EB53", x"EAF4", x"EADC",
		x"EAE4", x"EAFF", x"EB22", x"EB95", x"EC56", x"ED8C", x"EFA7", x"F362",
		x"F907", x"008B", x"0892", x"0F43", x"12E0", x"1333", x"1171", x"0F9D",
		x"0F2C", x"1064", x"120B", x"125D", x"0FBD", x"09EE", x"0245", x"FB57",
		x"F79A", x"F858", x"FD40", x"0494", x"0C0F", x"1177", x"1393", x"12AE",
		x"0FE4", x"0CF4", x"0B23", x"0AFB", x"0C47", x"0E7D", x"1124", x"138B",
		x"14D8", x"1453", x"1151", x"0BB9", x"0450", x"FC40", x"F4D7", x"EF5F",
		x"EC07", x"EAA8", x"EA69", x"EAD2", x"EB64", x"EC3F", x"ED9D", x"EF80",
		x"F14E", x"F2A0", x"F317", x"F2D1", x"F1D1", x"F062", x"EEB4", x"ECE7",
		x"EB8A", x"EAE1", x"EB06", x"EBBB", x"ECEF", x"EEB7", x"F0F3", x"F357",
		x"F50E", x"F580", x"F468", x"F1F8", x"EF22", x"ECF2", x"ECF5", x"EFDA",
		x"F58C", x"FCBE", x"0417", x"0A3A", x"0E9D", x"1136", x"1269", x"12F8",
		x"134D", x"13DF", x"1466", x"14BE", x"14C1", x"1415", x"12BA", x"10D7",
		x"0EC9", x"0D75", x"0D49", x"0EA0", x"10E9", x"1313", x"13EC", x"1288",
		x"0E75", x"0829", x"0099", x"F933", x"F31C", x"EEF0", x"EC70", x"EB27",
		x"EAA4", x"EA9F", x"EADC", x"EB0E", x"EB6D", x"EC76", x"EEC9", x"F2F2",
		x"F92A", x"00A0", x"086B", x"0EE3", x"1292", x"128E", x"0EAE", x"07E9",
		x"FFF7", x"F888", x"F296", x"EEAE", x"EC58", x"EB70", x"EB6B", x"EC41",
		x"EDE0", x"F023", x"F29D", x"F4C7", x"F5D0", x"F50A", x"F285", x"EF4E",
		x"ECED", x"ED2D", x"F0DB", x"F75A", x"FEBE", x"0593", x"0AAA", x"0DFA",
		x"0FE3", x"10C8", x"1158", x"11FE", x"1312", x"1448", x"148B", x"12C2",
		x"0E2D", x"0716", x"FECF", x"F70B", x"F112", x"ED55", x"EB99", x"EB28",
		x"EBA5", x"ECC2", x"EE50", x"F074", x"F2E8", x"F55A", x"F734", x"F82F",
		x"F7F8", x"F6BF", x"F4B1", x"F239", x"EF8E", x"ED4B", x"EBEA", x"EBC6",
		x"ED38", x"F06C", x"F565", x"FC04", x"0397", x"0AF9", x"10CC", x"13DB",
		x"1376", x"0FC5", x"0995", x"0229", x"FAE7", x"F48B", x"EF8D", x"EC51",
		x"EAD6", x"EACC", x"EB8A", x"EC6F", x"ED20", x"EDCD", x"EEA3", x"F010",
		x"F237", x"F542", x"F8FE", x"FD54", x"019A", x"0508", x"06A9", x"063A",
		x"035E", x"FE1A", x"F773", x"F0FA", x"ED1D", x"ED01", x"EFE6", x"F375",
		x"F588", x"F4F1", x"F213", x"EF0C", x"EE38", x"F111", x"F6D3", x"FD59",
		x"01C0", x"0212", x"FE15", x"F765", x"F12D", x"EDD2", x"EE68", x"F189",
		x"F4DE", x"F659", x"F500", x"F1A5", x"EE42", x"ED7B", x"F0A6", x"F6F0",
		x"FE05", x"0368", x"05D3", x"0543", x"0277", x"FE55", x"F9DB", x"F5EE",
		x"F313", x"F17D", x"F165", x"F2AC", x"F4E8", x"F7C7", x"FB1C", x"FE3F",
		x"00CB", x"0272", x"031C", x"02EF", x"01D3", x"FFC0", x"FCDD", x"F98B",
		x"F62F", x"F33B", x"F0E4", x"EF25", x"EDBB", x"EC83", x"EB77", x"EAC8",
		x"EAAB", x"EAE9", x"EB6C", x"EC70", x"EDED", x"EFE2", x"F237", x"F4B3",
		x"F6F1", x"F8BA", x"F9A6", x"F983", x"F845", x"F66B", x"F41A", x"F1CE",
		x"EF95", x"EDC7", x"ECA5", x"EC04", x"EBDA", x"EC17", x"ECBD", x"EDC5",
		x"EF6E", x"F1E9", x"F58B", x"FA62", x"002E", x"066A", x"0C6C", x"114B",
		x"13EF", x"13C1", x"1091", x"0ABE", x"0320", x"FAE3", x"F38A", x"EE59",
		x"EC22", x"ECE7", x"EFFC", x"F467", x"F932", x"FDD5", x"020A", x"05A8",
		x"08AF", x"0B17", x"0CFA", x"0E7D", x"0FBC", x"10D5", x"11D8", x"12C4",
		x"13AC", x"146A", x"14ED", x"152E", x"149B", x"1269", x"0DDE", x"06C7",
		x"FE48", x"F653", x"F039", x"EC84", x"EACA", x"EA50", x"EACD", x"ECA3",
		x"F066", x"F65D", x"FE58", x"06E1", x"0E14", x"1269", x"12D0", x"0F42",
		x"088F", x"001C", x"F7E2", x"F14D", x"ED06", x"EACA", x"EA2B", x"EB0C",
		x"ED8D", x"F237", x"F8F9", x"011C", x"093C", x"0F6E", x"1270", x"119E",
		x"0D34", x"0634", x"FE0D", x"F63E", x"F046", x"ECBA", x"EB8E", x"EBB2",
		x"EC21", x"EC24", x"EB9A", x"EB42", x"EB84", x"EC87", x"EDBF", x"EE97",
		x"EEC2", x"EE2D", x"ECFE", x"EBCC", x"EADD", x"EAC3", x"EB4A", x"EC60",
		x"EDB7", x"EF24", x"F0CB", x"F298", x"F4A8", x"F711", x"F9D8", x"FCC7",
		x"FFA6", x"024A", x"04AA", x"06EB", x"0912", x"0B2F", x"0D4D", x"0F38",
		x"110F", x"129A", x"13E6", x"14DF", x"1522", x"1496", x"13DE", x"1363",
		x"1393", x"1447", x"14FA", x"1549", x"1501", x"142B", x"1345", x"12CF",
		x"1315", x"13BB", x"143A", x"13C6", x"1162", x"0C68", x"04D8", x"FC27",
		x"F45B", x"EEBB", x"EC20", x"EC73", x"EF8D", x"F4C1", x"FB63", x"02A3",
		x"098A", x"0F50", x"12F4", x"1381", x"1101", x"0BC3", x"0508", x"FDC4",
		x"F71B", x"F1CA", x"EE38", x"EC2F", x"EB30", x"EABF", x"EABD", x"EB16",
		x"EBA9", x"EC90", x"EDBA", x"EF49", x"F1A2", x"F500", x"F920", x"FD22",
		x"FFCC", x"001E", x"FDDE", x"F965", x"F3DF", x"EF3C", x"ED20", x"EE5B",
		x"F23D", x"F6EC", x"FA59", x"FB37", x"F95A", x"F567", x"F0F1", x"EDA3",
		x"ED28", x"F06A", x"F72A", x"0021", x"0943", x"1020", x"1363", x"12CB",
		x"0F6E", x"0ADE", x"06F3", x"0551", x"06A8", x"0A5E", x"0F15", x"129F",
		x"130B", x"1016", x"0AD0", x"0555", x"0156", x"0020", x"018E", x"04C7",
		x"08F4", x"0D02", x"1046", x"124E", x"12DB", x"1208", x"0FD6", x"0C99",
		x"08E3", x"0537", x"028D", x"01A0", x"02EB", x"0671", x"0B3B", x"1007",
		x"12E8", x"12F0", x"0FEB", x"0ACE", x"04C0", x"FEE5", x"F9E4", x"F62E",
		x"F3A3", x"F1E2", x"F097", x"EF58", x"EE44", x"ED21", x"EC30", x"EB79",
		x"EB0C", x"EB3E", x"EBF1", x"ECE7", x"EDAB", x"EDEB", x"EDA4", x"ECE6",
		x"EC1B", x"EBB4", x"EBC2", x"EBFD", x"EC42", x"EC75", x"EC52", x"EBF1",
		x"EB81", x"EB3B", x"EB6A", x"EC08", x"ECB8", x"ECE7", x"EC8C", x"EC0D",
		x"EC23", x"EDA4", x"F147", x"F788", x"FF97", x"07F8", x"0EEC", x"12E2",
		x"132E", x"0FD4", x"09B6", x"0262", x"FB5E", x"F5E4", x"F20D", x"EFE5",
		x"EF17", x"EF79", x"F0CB", x"F34A", x"F6CC", x"FAED", x"FF2C", x"02D7",
		x"05F0", x"0873", x"0A8D", x"0C41", x"0DCA", x"0F6D", x"1132", x"12F8",
		x"1485", x"1564", x"156A", x"14AB", x"1361", x"1229", x"11BC", x"1252",
		x"136C", x"13F9", x"12D6", x"0F40", x"090D", x"011F", x"F91E", x"F2E7",
		x"EFA0", x"EF20", x"F0C5", x"F3B8", x"F7BA", x"FC0E", x"FFDB", x"01C6",
		x"0103", x"FD2F", x"F757", x"F186", x"EDEE", x"EDE2", x"F0D4", x"F4F9",
		x"F81C", x"F897", x"F647", x"F239", x"EE59", x"ECFC", x"EF03", x"F427",
		x"FAEC", x"01C1", x"079A", x"0BFE", x"0F14", x"110F", x"1241", x"12F3",
		x"133D", x"1322", x"12E9", x"1244", x"1151", x"0FD8", x"0DEB", x"0B41",
		x"07F7", x"048C", x"010F", x"FE12", x"FB7B", x"F959", x"F760", x"F5A4",
		x"F3D7", x"F1F2", x"F00F", x"EE02", x"EC3E", x"EB3E", x"EB0C", x"EB43",
		x"EB82", x"EB38", x"EAC1", x"EB0B", x"ECFD", x"F11D", x"F785", x"FF42",
		x"071E", x"0DB4", x"121A", x"1405", x"1412", x"12AB", x"1075", x"0DBA",
		x"0AC2", x"07F1", x"0654", x"06DD", x"0999", x"0DB1", x"1194", x"1373",
		x"1218", x"0D69", x"063B", x"FDEB", x"F5F6", x"EFBE", x"EC3B", x"EBE3",
		x"EE8D", x"F342", x"F908", x"FEF9", x"049D", x"0971", x"0D30", x"0FCF",
		x"116B", x"1259", x"12FB", x"135F", x"13A3", x"139A", x"12E4", x"117F",
		x"0F8B", x"0D2C", x"0AA6", x"07E9", x"0539", x"027A", x"0002", x"FE16",
		x"FCB1", x"FB46", x"F92B", x"F60F", x"F263", x"EEEF", x"ED28", x"EE25",
		x"F21E", x"F874", x"FFB3", x"0671", x"0B11", x"0C4E", x"0978", x"0356",
		x"FB92", x"F441", x"EF2B", x"ECD9", x"ECE5", x"EE3F", x"EFBA", x"EFFD",
		x"EEEB", x"ED35", x"EBAB", x"EAD1", x"EAA6", x"EAC4", x"EB1A", x"EBFA",
		x"EE3D", x"F25C", x"F8D0", x"00E3", x"0937", x"0FCE", x"1366", x"1348",
		x"0F78", x"0909", x"013F", x"F970", x"F30C", x"EEAE", x"EC7B", x"EBBD",
		x"EBF9", x"ECFB", x"EECB", x"F16F", x"F44D", x"F6E6", x"F88D", x"F90C",
		x"F840", x"F655", x"F3D0", x"F0FC", x"EE8F", x"ECC1", x"EBC2", x"EB90",
		x"EBB5", x"EC03", x"EC82", x"ED68", x"EF07", x"F180", x"F53D", x"FA44",
		x"006F", x"075E", x"0DD6", x"1254", x"13C2", x"1233", x"0E8F", x"0A9E",
		x"07EC", x"0747", x"08F7", x"0BFE", x"0F38", x"11DC", x"1394", x"1483",
		x"14BB", x"1463", x"13B3", x"126B", x"108F", x"0E47", x"0BEE", x"0A04",
		x"08C3", x"085D", x"0897", x"0983", x"0B1D", x"0D0C", x"0F09", x"111E",
		x"12E8", x"1386", x"11FE", x"0DB1", x"0704", x"FF36", x"F7BD", x"F19F",
		x"EDA2", x"EBB7", x"EB24", x"EB4E", x"EBD3", x"ECF0", x"EEC8", x"F145",
		x"F457", x"F7E5", x"FB9B", x"FF40", x"0280", x"0532", x"0767", x"0922",
		x"0A36", x"0ACA", x"0B2C", x"0B3E", x"0B0E", x"0A45", x"0871", x"0588",
		x"015D", x"FC16", x"F634", x"F0D1", x"ED2F", x"EC30", x"EE1B", x"F268",
		x"F818", x"FDE0", x"02BC", x"05F5", x"077D", x"077D", x"0601", x"034A",
		x"FF56", x"FA63", x"F526", x"F052", x"ECEA", x"EBF7", x"EDE8", x"F286",
		x"F8F0", x"FFA7", x"0589", x"09C5", x"0C28", x"0CD7", x"0C4D", x"0ABA",
		x"07ED", x"033D", x"FCBA", x"F602", x"F1E7", x"F258", x"F681", x"FAAF",
		x"FB51", x"F76B", x"F178", x"EC9B", x"EA66", x"EA53", x"EAF1", x"EB6F",
		x"EC27", x"EDAB", x"F064", x"F4B2", x"FA69", x"010B", x"07CA", x"0DD0",
		x"1217", x"13F7", x"130C", x"0FB9", x"0B15", x"065F", x"0270", x"FF95",
		x"FDD5", x"FC72", x"FAEB", x"F897", x"F547", x"F185", x"EE2D", x"EC98",
		x"ED92", x"F173", x"F7C2", x"FF15", x"060E", x"0B73", x"0EFC", x"1104",
		x"1248", x"1334", x"13EC", x"1463", x"14BA", x"1483", x"131B", x"0FE0",
		x"0A91", x"03B0", x"FC23", x"F50F", x"EF76", x"EC80", x"ECB1", x"F005",
		x"F58E", x"FC6D", x"0389", x"0A46", x"0FC2", x"1320", x"13D9", x"11CD",
		x"0D39", x"06BB", x"FF5D", x"F81D", x"F202", x"EDEA", x"EC33", x"ED0B",
		x"F07E", x"F62F", x"FD50", x"04E5", x"0BCE", x"1100", x"13A7", x"138B",
		x"1097", x"0B8A", x"0525", x"FE52", x"F791", x"F1BE", x"EDAD", x"EC94",
		x"EF24", x"F52B", x"FD49", x"05A7", x"0CC0", x"11A9", x"1481", x"158E",
		x"151D", x"1338", x"0F67", x"0960", x"0160", x"F8D3", x"F1B8", x"EDA0",
		x"ED1B", x"EFC9", x"F4F7", x"FBB5", x"02DB", x"0966", x"0ED4", x"127D",
		x"13CE", x"126C", x"0E57", x"0837", x"00F7", x"F99B", x"F30F", x"EE5D",
		x"EC20", x"ECB6", x"F017", x"F58D", x"FC7A", x"03BB", x"0A7F", x"0FF6",
		x"1339", x"1346", x"0F42", x"0800", x"FF17", x"F6C5", x"F087", x"ECB6",
		x"EAEA", x"EAD0", x"ECE4", x"F128", x"F779", x"FF48", x"0737", x"0E15",
		x"12EA", x"1542", x"1542", x"1357", x"0F7E", x"095E", x"012B", x"F84B",
		x"F0E4", x"ECEE", x"ECEC", x"F06B", x"F5F0", x"FC7F", x"0328", x"0979",
		x"0EFF", x"12AC", x"13AA", x"115C", x"0C2D", x"0503", x"FD2D", x"F605",
		x"F060", x"ECC1", x"EB47", x"EB51", x"EC32", x"ED99", x"EF2C", x"F114",
		x"F2FC", x"F4CD", x"F660", x"F7DA", x"F93B", x"FAC8", x"FCC3", x"FF68",
		x"02AF", x"064C", x"0A20", x"0DBC", x"10E6", x"132C", x"13C4", x"11DE",
		x"0D2C", x"0612", x"FDD7", x"F623", x"F014", x"EC86", x"EBDE", x"EDE0",
		x"F21F", x"F820", x"FF52", x"06C5", x"0D4B", x"1197", x"1266", x"0F9C",
		x"09B9", x"025C", x"FBB0", x"F792", x"F739", x"FAE1", x"0164", x"08E9",
		x"0F1B", x"1270", x"12C4", x"118E", x"105C", x"1033", x"1130", x"11E0",
		x"1037", x"0B21", x"0380", x"FBBC", x"F6A3", x"F638", x"FA87", x"0217",
		x"0A42", x"1052", x"131C", x"1309", x"11CB", x"110F", x"1156", x"12B1",
		x"1362", x"11C8", x"0CD0", x"0533", x"FCDA", x"F5B4", x"F0A2", x"EDAF",
		x"EC12", x"EB4E", x"EB01", x"EADA", x"EADB", x"EAEA", x"EB18", x"EBB3",
		x"ECB1", x"EE60", x"F05E", x"F250", x"F46C", x"F68E", x"F8F0", x"FB41",
		x"FDA2", x"0006", x"02A8", x"056C", x"0830", x"0AC7", x"0D16", x"0EF8",
		x"1072", x"119B", x"125D", x"132C", x"13ED", x"14B6", x"14D0", x"1307",
		x"0E7C", x"0723", x"FE58", x"F614", x"EFDE", x"EC28", x"EA83", x"EA39",
		x"EB75", x"EED2", x"F461", x"FBD7", x"040A", x"0BA7", x"1131", x"13FD",
		x"1401", x"119B", x"0D2C", x"06A2", x"FE4F", x"F5EC", x"EF5C", x"EC7D",
		x"EDA7", x"F208", x"F819", x"FECB", x"0567", x"0B92", x"107B", x"1340",
		x"132E", x"0FB2", x"0904", x"0056", x"F7B9", x"F0F2", x"ECEC", x"EAFB",
		x"EA65", x"EA4F", x"EA6F", x"EAB2", x"EB1E", x"EBCA", x"ECD2", x"EE43",
		x"EFC7", x"F0DA", x"F151", x"F0F6", x"EFDC", x"EE40", x"EC92", x"EB61",
		x"EB4D", x"ECCF", x"EFF5", x"F4C7", x"FAE0", x"01C3", x"08BF", x"0EAE",
		x"1280", x"132F", x"10A3", x"0B2E", x"03E9", x"FC42", x"F54E", x"EFE3",
		x"EC6C", x"EAE8", x"EB2B", x"ECEC", x"EF84", x"F26A", x"F505", x"F711",
		x"F85E", x"F8EA", x"F892", x"F726", x"F4B3", x"F1AE", x"EF04", x"ED14",
		x"EBFE", x"EB78", x"EC1B", x"EE8F", x"F398", x"FB01", x"035F", x"0AFD",
		x"10C4", x"146C", x"161E", x"1621", x"147A", x"10B8", x"0AD1", x"031C",
		x"FAA7", x"F2DF", x"ED72", x"EB89", x"ED75", x"F288", x"F9C2", x"01E1",
		x"0997", x"0FD9", x"13BD", x"1555", x"157E", x"1529", x"1503", x"14DA",
		x"1428", x"12C7", x"111F", x"0FEB", x"0F7A", x"1036", x"11B8", x"1331",
		x"1458", x"14E2", x"1504", x"14F3", x"14F4", x"14EF", x"14E7", x"14BC",
		x"1424", x"132E", x"1206", x"1109", x"104E", x"1028", x"107A", x"114D",
		x"1272", x"13B8", x"14C5", x"1533", x"14F3", x"13FF", x"1272", x"1081",
		x"0E31", x"0BB5", x"0942", x"074F", x"0660", x"067F", x"078B", x"0939",
		x"0B88", x"0E12", x"1070", x"1228", x"1332", x"13B1", x"13D1", x"1395",
		x"129E", x"10D6", x"0E51", x"0B48", x"0812", x"04F8", x"0232", x"FFF6",
		x"FE38", x"FCD0", x"FB53", x"F921", x"F63C", x"F2CF", x"EF7B", x"ED14",
		x"EC73", x"EE7F", x"F320", x"F9C0", x"0125", x"081C", x"0DA8", x"115D",
		x"136C", x"1465", x"14EE", x"153F", x"1533", x"14C6", x"1427", x"1364",
		x"12B2", x"11E5", x"10F0", x"0F76", x"0D44", x"0A00", x"05BB", x"009B",
		x"FB09", x"F565", x"F083", x"ED16", x"EC04", x"EDF7", x"F30E", x"FAB5",
		x"033B", x"0B17", x"10A3", x"1321", x"1270", x"0F8C", x"0BF1", x"094E",
		x"0904", x"0B0A", x"0E70", x"11D8", x"1381", x"121D", x"0D54", x"05A7",
		x"FC99", x"F41F", x"EE64", x"ECB8", x"EF09", x"F3EC", x"F946", x"FD4E",
		x"FE5E", x"FC4D", x"F781", x"F205", x"EE2B", x"ED9C", x"F044", x"F48D",
		x"F7F7", x"F8BD", x"F682", x"F263", x"EE8E", x"ED63", x"EFB7", x"F4E4",
		x"FAF2", x"0003", x"02FC", x"03B0", x"0231", x"FF41", x"FB53", x"F704",
		x"F298", x"EEC9", x"EC41", x"EBB7", x"EDAA", x"F23A", x"F8F1", x"0088",
		x"07DD", x"0DA9", x"11B3", x"13DB", x"14CA", x"1500", x"1503", x"14EC",
		x"14BB", x"142F", x"1331", x"1205", x"10CA", x"0F64", x"0D9E", x"0B69",
		x"08B0", x"05A1", x"024B", x"FEE5", x"FB7B", x"F810", x"F4D0", x"F231",
		x"F05D", x"EFA6", x"F01D", x"F24A", x"F617", x"FB9E", x"0256", x"094D",
		x"0F35", x"129E", x"12AC", x"0F45", x"0969", x"024F", x"FB40", x"F4F2",
		x"F005", x"ED05", x"EC70", x"EEC8", x"F44B", x"FC8E", x"05E1", x"0DF3",
		x"1300", x"14AF", x"1495", x"142C", x"145A", x"148C", x"13D1", x"1143",
		x"0C44", x"0526", x"FCEE", x"F54D", x"EFA2", x"EC75", x"EB7B", x"EBE8",
		x"ECD6", x"EDC3", x"EDDD", x"ED18", x"EBC3", x"EB1F", x"EC4F", x"F003",
		x"F622", x"FDAB", x"057B", x"0C07", x"1015", x"10CF", x"0E2F", x"08D3",
		x"01CD", x"FA14", x"F30B", x"EE19", x"EC43", x"ED4D", x"F017", x"F2C7",
		x"F476", x"F52B", x"F5A9", x"F717", x"FA15", x"FEFD", x"052A", x"0B99",
		x"10BD", x"135D", x"12B2", x"0F3A", x"0A84", x"0630", x"035C", x"027A",
		x"0304", x"04BD", x"0771", x"0A89", x"0D91", x"1014", x"1238", x"13AE",
		x"147F", x"1463", x"13BA", x"12C6", x"1210", x"122F", x"1319", x"13E6",
		x"135F", x"104A", x"0A9A", x"032C", x"FB63", x"F4CA", x"F08E", x"EFBF",
		x"F267", x"F814", x"FFA1", x"078B", x"0E50", x"128A", x"139C", x"122A",
		x"0F74", x"0CC6", x"0B02", x"0A08", x"0922", x"077F", x"0493", x"0010",
		x"FA79", x"F48A", x"EFAC", x"ED53", x"EDF4", x"F160", x"F634", x"FACF",
		x"FD9D", x"FE56", x"FCCB", x"F9E4", x"F63D", x"F2B7", x"F001", x"EE6B",
		x"EDC3", x"EE4F", x"F00E", x"F2F1", x"F6DD", x"FAEF", x"FDF4", x"FF09",
		x"FD89", x"F9B9", x"F493", x"EFD1", x"ED5A", x"EE30", x"F22A", x"F76F",
		x"FB68", x"FC48", x"F99E", x"F4D7", x"F03C", x"EDB7", x"EE63", x"F252",
		x"F85A", x"FEC9", x"0444", x"083E", x"0ACC", x"0C87", x"0D9B", x"0E9E",
		x"0FCF", x"1143", x"12C1", x"1410", x"14E8", x"1525", x"1506", x"14A1",
		x"1419", x"13CA", x"1399", x"13D8", x"1477", x"14F4", x"14CA", x"13F5",
		x"12F2", x"124C", x"124A", x"12E0", x"13DB", x"14B6", x"14C9", x"143A",
		x"1381", x"137B", x"1409", x"1430", x"12BD", x"0EEE", x"08CC", x"010D",
		x"F903", x"F282", x"EEA2", x"EE72", x"F1D9", x"F80E", x"FFE6", x"07E1",
		x"0EA6", x"1322", x"1506", x"14F2", x"1406", x"137D", x"139B", x"1429",
		x"1471", x"140E", x"12CC", x"10CA", x"0EBE", x"0CEB", x"0B4A", x"09AE",
		x"07B0", x"0553", x"029C", x"FFA1", x"FC67", x"F946", x"F637", x"F372",
		x"F0F3", x"EEF7", x"EDDB", x"ED6F", x"ED7C", x"EDF0", x"EF05", x"F0C6",
		x"F347", x"F64E", x"F956", x"FB9C", x"FC87", x"FBA8", x"F94C", x"F607",
		x"F2A6", x"EFB1", x"ED5C", x"EC13", x"EC3A", x"EEB1", x"F3BE", x"FB29",
		x"0387", x"0B14", x"10A3", x"13F8", x"1574", x"15F9", x"158F", x"1400",
		x"1094", x"0AD5", x"0307", x"FA80", x"F2FC", x"EDE0", x"EB66", x"EAC9",
		x"EB0F", x"EBB3", x"EC54", x"ECE5", x"ED77", x"EE33", x"EF79", x"F156",
		x"F3C3", x"F689", x"F950", x"FBF9", x"FE76", x"00DE", x"0391", x"0674",
		x"0973", x"0C6B", x"0F25", x"114D", x"12B3", x"1368", x"1386", x"12E8",
		x"116B", x"0EF2", x"0BBA", x"0876", x"05BD", x"046C", x"0508", x"07C8",
		x"0C18", x"1021", x"1228", x"10D2", x"0C56", x"066B", x"01A5", x"000E",
		x"0287", x"0807", x"0E1A", x"122A", x"1269", x"0F7A", x"0B60", x"089A",
		x"08B6", x"0BAD", x"0FC7", x"12A3", x"125D", x"0E53", x"07AB", x"008A",
		x"FA5F", x"F5E4", x"F2F5", x"F10C", x"EFED", x"EF19", x"EE3B", x"ED02",
		x"EBDE", x"EB0B", x"EAD6", x"EB4B", x"EC40", x"ED74", x"EE96", x"EF43",
		x"EF48", x"EEC1", x"EDCC", x"ECD3", x"EBF1", x"EB57", x"EB19", x"EB1D",
		x"EB12", x"EB18", x"EB06", x"EAE9", x"EAC3", x"EAB3", x"EAFB", x"EC08",
		x"EE77", x"F30D", x"F9C6", x"01E3", x"09EC", x"1030", x"1366", x"13ED",
		x"1314", x"1270", x"12A1", x"1355", x"1327", x"10B8", x"0B48", x"039F",
		x"FB94", x"F53C", x"F199", x"F056", x"F123", x"F37D", x"F707", x"FB4E",
		x"FFD4", x"0410", x"0769", x"09CC", x"0B59", x"0C78", x"0D92", x"0EDE",
		x"108C", x"1272", x"13DE", x"13B9", x"112E", x"0C1D", x"0554", x"FDC9",
		x"F698", x"F0E6", x"ED4C", x"EB94", x"EB4B", x"EC2C", x"EDAD", x"EFDD",
		x"F2AB", x"F597", x"F7D2", x"F8DB", x"F823", x"F5DB", x"F2C4", x"EF99",
		x"ED0A", x"EB50", x"EA72", x"EAD0", x"ED6B", x"F2CE", x"FABA", x"038E",
		x"0B64", x"111D", x"1481", x"1616", x"1615", x"1477", x"10F9", x"0B72",
		x"0404", x"FBB8", x"F3E3", x"EE3F", x"EB4F", x"EAC0", x"EB43", x"EC36",
		x"ED77", x"EF3C", x"F1CE", x"F4E9", x"F84F", x"FBC4", x"FF39", x"02B1",
		x"05AF", x"082A", x"0A17", x"0B93", x"0C69", x"0C57", x"0B40", x"0940",
		x"0676", x"0344", x"FFDC", x"FCD7", x"FABF", x"F9F0", x"FA84", x"FC89",
		x"FF79", x"02FC", x"06A6", x"09F8", x"0C2B", x"0CFD", x"0C1E", x"09BD",
		x"0616", x"020D", x"FE2A", x"FB06", x"F963", x"F9D0", x"FCAC", x"020C",
		x"08B8", x"0EDC", x"12A9", x"1340", x"10FD", x"0D75", x"0A35", x"083F",
		x"0815", x"09A5", x"0C78", x"0FA6", x"1245", x"140C", x"14C9", x"14F5",
		x"14BB", x"1456", x"13C7", x"12CA", x"1166", x"0FAB", x"0DB9", x"0B6B",
		x"090A", x"069D", x"044F", x"0231", x"FFE5", x"FD69", x"FA9B", x"F7A3",
		x"F4AD", x"F20F", x"EFBE", x"EDDB", x"EC6E", x"EBA1", x"EB5F", x"EB5C",
		x"EB71", x"EB8E", x"EBB2", x"EBFB", x"EC8A", x"EE18", x"F11B", x"F60A",
		x"FC7B", x"03DF", x"0B34", x"10F2", x"13D5", x"138F", x"1104", x"0E45",
		x"0CED", x"0DB8", x"0FFB", x"125D", x"12FC", x"109A", x"0AE5", x"02EE",
		x"FA4C", x"F2C6", x"EDC2", x"EC0D", x"EDAB", x"F1D9", x"F7A3", x"FDED",
		x"03EA", x"08DC", x"0C89", x"0EF1", x"1056", x"114C", x"124B", x"1372",
		x"1488", x"14A6", x"12DC", x"0E7B", x"07C3", x"FFA9", x"F79C", x"F0DE",
		x"EC85", x"EA94", x"EA76", x"EB2E", x"EC84", x"EE3A", x"F04D", x"F25A",
		x"F3DA", x"F415", x"F2CB", x"F065", x"EDB2", x"EC3A", x"ED31", x"F145",
		x"F82D", x"00D8", x"0981", x"100F", x"12F9", x"11E7", x"0D84", x"076E",
		x"014C", x"FCCB", x"FAD5", x"FC2D", x"0078", x"06B2", x"0CF0", x"1181",
		x"12FB", x"115D", x"0D73", x"0870", x"0384", x"FF88", x"FCD1", x"FAF8",
		x"F990", x"F808", x"F662", x"F499", x"F321", x"F1D8", x"F083", x"EF20",
		x"ED9F", x"EC41", x"EB27", x"EB0A", x"EC8A", x"F06F", x"F6D6", x"FEB7",
		x"06BE", x"0D58", x"11F1", x"1471", x"155B", x"1547", x"14DF", x"1489",
		x"143D", x"1376", x"11A4", x"0E0A", x"086F", x"010C", x"F8D5", x"F195",
		x"ED42", x"EC79", x"EE23", x"F05B", x"F146", x"F082", x"EE9C", x"ED67",
		x"EE85", x"F2C4", x"F988", x"00B9", x"05A9", x"069A", x"0347", x"FCE1",
		x"F5A0", x"EFD7", x"ED29", x"EDA7", x"F050", x"F369", x"F5AB", x"F67C",
		x"F588", x"F34D", x"F06B", x"EDB6", x"EBE9", x"EB75", x"ECE2", x"F041",
		x"F578", x"FC29", x"0395", x"0A9D", x"1029", x"139A", x"14BA", x"1419",
		x"128C", x"10EE", x"0F77", x"0E36", x"0D62", x"0D04", x"0D58", x"0E0A",
		x"0EF2", x"0FE5", x"10F6", x"1223", x"1355", x"143F", x"14AC", x"1437",
		x"12F3", x"10FA", x"0EB6", x"0CB5", x"0B3C", x"0AEE", x"0BBF", x"0DB4",
		x"103E", x"129D", x"13AD", x"126B", x"0E3A", x"0743", x"FEB5", x"F638",
		x"EF84", x"EBEF", x"EBE5", x"EEBC", x"F350", x"F8E3", x"FEBE", x"0497",
		x"0A03", x"0E94", x"11F6", x"1426", x"1533", x"155A", x"1531", x"14A7",
		x"1334", x"1056", x"0BA5", x"0553", x"FDE5", x"F684", x"F071", x"ECB7",
		x"EB9E", x"ECA8", x"EEF9", x"F1DE", x"F4DF", x"F77C", x"F8CE", x"F82B",
		x"F5BA", x"F228", x"EEC4", x"ED28", x"EE92", x"F2E1", x"F92B", x"FF63",
		x"0388", x"0434", x"00E7", x"FABB", x"F3E2", x"EEB1", x"ECC5", x"EDFF",
		x"F14F", x"F519", x"F7DE", x"F8D7", x"F7DD", x"F58A", x"F25B", x"EF34",
		x"EC99", x"EB36", x"EBC7", x"EE9E", x"F3A0", x"FA4E", x"01D7", x"091F",
		x"0F12", x"130E", x"14C4", x"14D7", x"141D", x"1355", x"12AB", x"11D4",
		x"10B4", x"0F33", x"0D54", x"0AF3", x"07D2", x"03CE", x"FFAA", x"FC4D",
		x"FA1C", x"F92A", x"F952", x"FA55", x"FC6F", x"FFA2", x"035A", x"06F2",
		x"09C2", x"0B3D", x"0B46", x"0963", x"055C", x"FF6F", x"F8A5", x"F262",
		x"EE18", x"ECFC", x"EF97", x"F544", x"FC7B", x"03C2", x"0A2C", x"0F45",
		x"12D5", x"144C", x"1302", x"0EB9", x"07DF", x"FF9D", x"F75C", x"F0C2",
		x"ECBB", x"EB86", x"EC87", x"EE70", x"F039", x"F0EE", x"F06B", x"EF1C",
		x"ED8C", x"EC50", x"EB83", x"EB3B", x"EB8E", x"ECAB", x"EE8B", x"F158",
		x"F48E", x"F78E", x"F971", x"F95A", x"F757", x"F3B8", x"EFBD", x"ED44",
		x"EDAB", x"F142", x"F717", x"FD1D", x"0165", x"0235", x"FF88", x"FA32",
		x"F40E", x"EF50", x"ED65", x"EED5", x"F31C", x"F90A", x"FF54", x"04BC",
		x"08C2", x"0B6C", x"0D08", x"0DBF", x"0D9C", x"0BFD", x"0851", x"0269",
		x"FB35", x"F42B", x"EF15", x"EC9B", x"ECC5", x"EE86", x"F067", x"F12D",
		x"F05D", x"EE74", x"EC85", x"EB43", x"EAC8", x"EB0F", x"EB4B", x"EB42",
		x"EB10", x"EB75", x"ECCC", x"EEE0", x"F0C2", x"F15B", x"F059", x"EE5D",
		x"ECDF", x"ED31", x"F03E", x"F61C", x"FD7E", x"04C7", x"0A64", x"0DBD",
		x"0F0F", x"0E8C", x"0CA1", x"096D", x"0589", x"0150", x"FD46", x"F990",
		x"F640", x"F3B0", x"F1CA", x"F073", x"EF87", x"EE69", x"ED20", x"EBE3",
		x"EB2B", x"EB04", x"EB82", x"EC69", x"ED52", x"EE48", x"EEED", x"EF30",
		x"EEED", x"EE1D", x"ED0A", x"EC23", x"EB70", x"EB20", x"EB05", x"EB00",
		x"EB00", x"EADE", x"EA93", x"EA56", x"EA40", x"EA76", x"EB54", x"ED67",
		x"F146", x"F73D", x"FEC8", x"06D0", x"0DAF", x"1253", x"143D", x"1429",
		x"134F", x"1303", x"137A", x"13DC", x"1272", x"0E05", x"06C4", x"FE3A",
		x"F65A", x"F058", x"ECC1", x"EB23", x"EAD4", x"EAFC", x"EB29", x"EB57",
		x"EB84", x"EBC4", x"EC4A", x"ED35", x"EE84", x"F000", x"F19F", x"F3AA",
		x"F6BA", x"FAEE", x"0050", x"0685", x"0CAF", x"116A", x"1340", x"11C0",
		x"0DE5", x"0960", x"0626", x"0514", x"0669", x"096B", x"0D0A", x"1031",
		x"127E", x"13C5", x"1367", x"10CA", x"0B15", x"0336", x"FAA5", x"F34A",
		x"EE56", x"EB86", x"EA3E", x"EA15", x"EB71", x"EEB7", x"F433", x"FBCC",
		x"0437", x"0BD6", x"10F9", x"1297", x"1084", x"0B29", x"03D3", x"FBB7",
		x"F463", x"EF0B", x"EC16", x"EB51", x"EBAC", x"EC35", x"EC25", x"EB8B",
		x"EB37", x"EB5E", x"EC6D", x"EE44", x"F07C", x"F2C3", x"F4C1", x"F687",
		x"F83B", x"FA38", x"FCC0", x"FF93", x"028C", x"05AD", x"0913", x"0C3D",
		x"0EE1", x"10B4", x"11CE", x"1287", x"12EA", x"12BC", x"1204", x"10C0",
		x"0EFF", x"0CEA", x"0A99", x"07F7", x"04C4", x"00E0", x"FC8D", x"F84B",
		x"F4A7", x"F1C7", x"EFBE", x"EE95", x"EEBB", x"F0EA", x"F5B7", x"FCC8",
		x"04EA", x"0C39", x"114E", x"13C3", x"142D", x"13BD", x"1372", x"1365",
		x"12B7", x"0FDD", x"0A03", x"01B5", x"F90F", x"F1D5", x"ED43", x"EB15",
		x"EA8A", x"EA9B", x"EAD3", x"EADE", x"EB30", x"EC2D", x"EE92", x"F2C6",
		x"F8D3", x"004C", x"07E5", x"0E53", x"1295", x"146C", x"1408", x"11FB",
		x"0F10", x"0BC0", x"0887", x"059D", x"0349", x"01FC", x"01E3", x"030F",
		x"055F", x"0881", x"0BF8", x"0F1C", x"115E", x"1282", x"1275", x"10D2",
		x"0CE0", x"065A", x"FE25", x"F62E", x"EFF6", x"EC4B", x"EAE9", x"EAA3",
		x"EA9D", x"EAB3", x"EBD9", x"EF12", x"F523", x"FDA5", x"06B7", x"0E31",
		x"1290", x"1348", x"10B2", x"0B75", x"04AD", x"FD7E", x"F6FE", x"F1E0",
		x"EE61", x"EC32", x"EB33", x"EB10", x"EB84", x"EC44", x"ECE4", x"ED29",
		x"ECE9", x"EC72", x"EBAF", x"EAE9", x"EA8A", x"EAB1", x"EB5D", x"EBFD",
		x"EC51", x"EC06", x"EB82", x"EAEA", x"EAA1", x"EADA", x"EB83", x"EC3A",
		x"ECA8", x"EC43", x"EBC2", x"EBE4", x"EDBD", x"F1EF", x"F881", x"00A3",
		x"08E7", x"0F98", x"1305", x"1275", x"0E71", x"0803", x"00D0", x"F9F9",
		x"F48B", x"F0DC", x"EEF2", x"EE9D", x"EF8E", x"F1A4", x"F469", x"F79C",
		x"FA94", x"FD10", x"FE84", x"FEBC", x"FD9F", x"FB81", x"F8E0", x"F603",
		x"F334", x"F0A1", x"EE52", x"EC7F", x"EB50", x"EB02", x"EB5E", x"EC04",
		x"ECA0", x"ECCD", x"EC7A", x"EBF0", x"EBDB", x"ED66", x"F15C", x"F7C8",
		x"FFBF", x"077A", x"0D61", x"1099", x"1191", x"10B8", x"0E90", x"0B5E",
		x"0752", x"0374", x"0074", x"FF31", x"FFCA", x"0208", x"0562", x"0955",
		x"0CFB", x"0FB2", x"1106", x"10CE", x"0E8D", x"09FC", x"0395", x"FC2F",
		x"F4F0", x"EF44", x"EC1B", x"EBA2", x"EDAA", x"F14E", x"F54C", x"F907",
		x"FBBB", x"FD91", x"FED0", x"FF99", x"FFB5", x"FF03", x"FD90", x"FB9B",
		x"F975", x"F736", x"F4F7", x"F2B6", x"F073", x"EE4C", x"EC88", x"EB70",
		x"EB15", x"EB54", x"EBB3", x"EC04", x"EC37", x"EC0C", x"EBC1", x"EB78",
		x"EB69", x"EBBC", x"EC72", x"ED0B", x"ED2B", x"ECAD", x"EBF8", x"EBC6",
		x"ED22", x"F0B2", x"F689", x"FDF6", x"05AF", x"0C4B", x"1136", x"13E7",
		x"14DD", x"14B4", x"1419", x"139F", x"1395", x"140C", x"14A3", x"14D6",
		x"1379", x"0FD2", x"09BF", x"0207", x"FA17", x"F334", x"EE3B", x"EB5C",
		x"EA3A", x"EA3D", x"EAB6", x"EB72", x"EC1D", x"ECE7", x"EDF4", x"EFA9",
		x"F23D", x"F5B5", x"F9C0", x"FDB0", x"00A8", x"022D", x"01BE", x"FF4A",
		x"FAFC", x"F581", x"F063", x"ED3C", x"ED21", x"F000", x"F505", x"FABA",
		x"FFC7", x"037C", x"05AB", x"0711", x"0849", x"0A09", x"0C9E", x"0FAD",
		x"1261", x"140D", x"13DE", x"116C", x"0CB6", x"0613", x"FE37", x"F689",
		x"F052", x"ECEA", x"ED19", x"F0B0", x"F6C3", x"FE14", x"052E", x"0ABD",
		x"0E0F", x"0F10", x"0E20", x"0BE1", x"08A3", x"0510", x"01B8", x"FF69",
		x"FEBF", x"0045", x"0419", x"098B", x"0F34", x"12C9", x"1316", x"0FC0",
		x"0998", x"01E5", x"FA26", x"F366", x"EE68", x"EB78", x"EB13", x"ED55",
		x"F277", x"F9F2", x"0278", x"0A8D", x"107E", x"1340", x"12E4", x"1002",
		x"0C0E", x"08A6", x"06AC", x"0681", x"07DD", x"0A45", x"0CFC", x"0F90",
		x"1193", x"1301", x"13D1", x"1434", x"140B", x"137F", x"1258", x"106A",
		x"0D7F", x"0967", x"03D3", x"FD1C", x"F600", x"EFFD", x"ECB1", x"ECDA",
		x"EFC8", x"F3B5", x"F669", x"F69D", x"F464", x"F0E5", x"EE14", x"ED84",
		x"F026", x"F597", x"FCB1", x"03D5", x"09B9", x"0DD7", x"1050", x"11BB",
		x"12B8", x"1360", x"13DF", x"13E9", x"1380", x"1268", x"1075", x"0DB2",
		x"0AAC", x"07F4", x"0656", x"069C", x"08D1", x"0C4A", x"1010", x"1260",
		x"11A2", x"0D74", x"0734", x"00FA", x"FCB4", x"FB87", x"FD32", x"00C4",
		x"0534", x"0997", x"0CCC", x"0E55", x"0DB3", x"0A5F", x"0472", x"FCB3",
		x"F514", x"EF53", x"EC9B", x"EC8B", x"EE0F", x"EF92", x"F013", x"EF5D",
		x"EDF1", x"EC46", x"EB13", x"EA96", x"EABD", x"EB0A", x"EB33", x"EB1A",
		x"EB0F", x"EB9D", x"EC99", x"EE01", x"EF26", x"EFC9", x"EFC9", x"EF3D",
		x"EE49", x"ED22", x"EBFF", x"EB2F", x"EAA4", x"EAA8", x"EB34", x"EC4D",
		x"EDAF", x"EF36", x"F0C2", x"F27A", x"F4C3", x"F768", x"FA1D", x"FCB2",
		x"FF38", x"019C", x"0424", x"066A", x"08A7", x"0AFC", x"0D38", x"0F8B",
		x"11A6", x"1373", x"14A3", x"1518", x"1510", x"14D4", x"14BF", x"14C7",
		x"14E7", x"14FC", x"14D9", x"1471", x"1376", x"11D6", x"0F3C", x"0B4C",
		x"05E7", x"FF48", x"F826", x"F1B4", x"ED4B", x"EBB1", x"ED68", x"F1F7",
		x"F884", x"0018", x"075B", x"0D99", x"120C", x"142B", x"136F", x"0FFF",
		x"0A33", x"02A0", x"FA8D", x"F366", x"EE57", x"EBEE", x"EC2D", x"EE5B",
		x"F1B3", x"F522", x"F7E5", x"F9CA", x"FB1E", x"FC87", x"FEBD", x"024C",
		x"06D9", x"0BAD", x"0F9F", x"1149", x"0FC8", x"0B36", x"04F6", x"FF1E",
		x"FBED", x"FCA4", x"012B", x"07D3", x"0E5D", x"1286", x"1320", x"1119",
		x"0E38", x"0C5E", x"0CB5", x"0F25", x"122F", x"13A3", x"11B9", x"0BF7",
		x"039B", x"FA87", x"F2C8", x"EE0B", x"ED1C", x"EFB6", x"F4D4", x"FAB2",
		x"FFDC", x"02F6", x"031B", x"FFEB", x"FA73", x"F42E", x"EF18", x"ECA2",
		x"ED93", x"F164", x"F71C", x"FD06", x"01E6", x"055D", x"0774", x"08C2",
		x"0997", x"09D8", x"09EF", x"09C5", x"095D", x"08A5", x"0777", x"056B",
		x"0226", x"FDD4", x"F8A7", x"F35D", x"EF02", x"EC82", x"EC99", x"EF68",
		x"F48B", x"FB04", x"01AD", x"0759", x"0BCB", x"0EDC", x"10D8", x"11E7",
		x"12A2", x"135B", x"145B", x"14EE", x"13DB", x"104E", x"0A33", x"0267",
		x"FA35", x"F31E", x"EE17", x"EB4C", x"EA5E", x"EAD2", x"EBEE", x"EDD5",
		x"F031", x"F2E7", x"F4FB", x"F577", x"F40F", x"F13E", x"EE96", x"EDAB",
		x"EFAA", x"F4B4", x"FB6B", x"01A4", x"052C", x"04F5", x"014E", x"FB4A",
		x"F4CE", x"EF7C", x"ECEF", x"EE27", x"F2E5", x"FA4A", x"02CA", x"0AAD",
		x"108B", x"13B3", x"13ED", x"11E3", x"0E76", x"0A41", x"0603", x"0256",
		x"FF50", x"FCCD", x"FAAB", x"F8E0", x"F736", x"F57E", x"F3BC", x"F1FA",
		x"F04F", x"EED6", x"ED7F", x"EC5E", x"EB9A", x"EB38", x"EB3B", x"EBD7",
		x"ED2B", x"EF2C", x"F165", x"F352", x"F44E", x"F3FB", x"F263", x"EFF9",
		x"ED7D", x"EC04", x"EC89", x"EFFF", x"F666", x"FEDA", x"0797", x"0E8C",
		x"1239", x"11DE", x"0E00", x"07D2", x"00F8", x"FB52", x"F86A", x"F96B",
		x"FE42", x"0577", x"0CB5", x"11A0", x"135E", x"123C", x"1001", x"0E75",
		x"0EAD", x"1063", x"11F5", x"1198", x"0E1C", x"079D", x"FFA4", x"F7EE",
		x"F1D5", x"EDDD", x"EBE1", x"EB2E", x"EAE1", x"EA8A", x"EA3B", x"EA4D",
		x"EB49", x"EDEB", x"F284", x"F8E8", x"00A2", x"0854", x"0EAD", x"12F6",
		x"14FF", x"1562", x"151B", x"1476", x"135E", x"11A8", x"0F20", x"0BFA",
		x"08EC", x"060D", x"0406", x"0294", x"0178", x"FFEE", x"FD7F", x"F9DC",
		x"F56D", x"F0D2", x"ED58", x"EC24", x"EDDF", x"F253", x"F899", x"FF3A",
		x"04F8", x"08F4", x"0AD3", x"0AD5", x"094D", x"06A9", x"02DF", x"FE87",
		x"FA3A", x"F68E", x"F3F5", x"F238", x"F123", x"F048", x"EF80", x"EE76",
		x"ED17", x"EBF6", x"EC2F", x"EF16", x"F527", x"FD66", x"0609", x"0D3C",
		x"1239", x"14B7", x"14F0", x"12BC", x"0E60", x"0813", x"0060", x"F856",
		x"F157", x"ECB0", x"EAAF", x"EA74", x"EAD8", x"EB2A", x"EB3A", x"EB85",
		x"EC87", x"EEA8", x"F26E", x"F850", x"FFF9", x"07F5", x"0EB9", x"12BF",
		x"13E9", x"12D7", x"114E", x"10A3", x"115B", x"12DC", x"1358", x"1108",
		x"0B27", x"0313", x"FB11", x"F52B", x"F258", x"F271", x"F4C6", x"F8A7",
		x"FD4D", x"01CF", x"054C", x"0737", x"0728", x"054B", x"01ED", x"FDCC",
		x"F997", x"F634", x"F417", x"F3C7", x"F592", x"F9BB", x"FFC3", x"06D1",
		x"0D6B", x"1206", x"13AC", x"1264", x"0EE3", x"0A44", x"059C", x"01A1",
		x"FEA3", x"FC68", x"FADC", x"F9EA", x"F998", x"FA33", x"FBC5", x"FE1C",
		x"0108", x"043A", x"0778", x"0A38", x"0C14", x"0CB7", x"0BEA", x"0A00",
		x"071A", x"038C", x"FFBE", x"FC5C", x"FA0B", x"F960", x"FA40", x"FCDE",
		x"006B", x"046D", x"0817", x"0ACB", x"0C57", x"0C27", x"09C5", x"0517",
		x"FEAE", x"F789", x"F15C", x"ED90", x"EC91", x"EE3B", x"F1AB", x"F5FA",
		x"FA33", x"FDDC", x"008B", x"0257", x"0388", x"041F", x"0446", x"03E8",
		x"02D4", x"0109", x"FEA9", x"FBE6", x"F8C9", x"F5DB", x"F2F4", x"F066",
		x"EE8E", x"ED29", x"EC4C", x"EBB5", x"EB58", x"EB22", x"EB1C", x"EB6C",
		x"EC80", x"EEAA", x"F19C", x"F4C8", x"F767", x"F8D2", x"F8A3", x"F6DF",
		x"F3D9", x"F037", x"ED28", x"EC17", x"EDE0", x"F265", x"F8E3", x"0006",
		x"06B6", x"0C25", x"100C", x"1260", x"1353", x"139F", x"1396", x"1350",
		x"127D", x"1051", x"0C70", x"069E", x"FF71", x"F7D3", x"F150", x"ED51",
		x"ECC1", x"EFDD", x"F5D8", x"FD3E", x"04BA", x"0B34", x"1016", x"1336",
		x"1469", x"13D3", x"119F", x"0E9F", x"0B47", x"0845", x"0616", x"0576",
		x"066A", x"08F3", x"0C7B", x"103C", x"12EE", x"1335", x"1085", x"0B19",
		x"0474", x"FDB5", x"F822", x"F42D", x"F20B", x"F151", x"F0E5", x"EFF6",
		x"EE34", x"EC5A", x"EB82", x"ED08", x"F168", x"F858", x"008A", x"0857",
		x"0E70", x"1203", x"1297", x"1050", x"0B88", x"04E4", x"FD25", x"F59F",
		x"EF9A", x"EBFF", x"EAE1", x"EB41", x"EBE9", x"EBF7", x"EB75", x"EB00",
		x"EB84", x"ED51", x"F04F", x"F46F", x"F9C0", x"001D", x"06E1", x"0D27",
		x"11AF", x"139A", x"1256", x"0DF7", x"0725", x"FF0E", x"F742", x"F0F4",
		x"ECE8", x"EB49", x"EBD8", x"EE16", x"F13E", x"F4F0", x"F8BD", x"FC91",
		x"FFFA", x"024F", x"0359", x"030B", x"01B0", x"FF15", x"FBC2", x"F81B",
		x"F4E1", x"F29D", x"F158", x"F119", x"F255", x"F544", x"F9FA", x"0031",
		x"073A", x"0DF7", x"12AA", x"13C8", x"1081", x"0995", x"0090", x"F7B2",
		x"F0CF", x"ECBA", x"EB54", x"EB75", x"EBD6", x"EBCF", x"EBB3", x"EC62",
		x"EEF1", x"F431", x"FBB3", x"0408", x"0B1B", x"0F89", x"10F3", x"1024",
		x"0DE7", x"0A85", x"0677", x"023A", x"FEC8", x"FD0D", x"FD80", x"0017",
		x"0434", x"08BF", x"0CA4", x"0F49", x"107A", x"0FF0", x"0D20", x"07E2",
		x"00CF", x"F919", x"F23B", x"EDAB", x"EB86", x"EB6C", x"EC75", x"ED95",
		x"EE15", x"EDB5", x"EC90", x"EB6E", x"EAF2", x"EB61", x"EC92", x"EE6C",
		x"F0AA", x"F309", x"F56B", x"F7B8", x"F9B6", x"FB2F", x"FBCB", x"FB4D",
		x"F9FD", x"F7D6", x"F526", x"F264", x"F012", x"EE72", x"ED96", x"ED6E",
		x"EE14", x"EF42", x"F0F5", x"F34A", x"F60B", x"F8B9", x"FADD", x"FC1A",
		x"FC63", x"FBDA", x"FAA1", x"F8EA", x"F6E2", x"F45C", x"F160", x"EE56",
		x"EC40", x"EC28", x"EEBE", x"F408", x"FB32", x"0300", x"09F6", x"0EF2",
		x"11BC", x"1285", x"1214", x"10A3", x"0E5D", x"0B5D", x"07D8", x"0467",
		x"0119", x"FE0B", x"FB36", x"F89B", x"F656", x"F42D", x"F22E", x"F045",
		x"EEBB", x"ED80", x"EC97", x"EBD0", x"EB47", x"EAE0", x"EABE", x"EAF5",
		x"EC15", x"EED6", x"F3BD", x"FAD3", x"02E8", x"0A8C", x"1054", x"13C0",
		x"14DD", x"1463", x"132E", x"1274", x"1263", x"1323", x"140F", x"14AC",
		x"145F", x"1274", x"0E53", x"07BB", x"FF83", x"F70D", x"F076", x"EC6E",
		x"EADB", x"EAC1", x"EB13", x"EB2D", x"EB6B", x"ECC3", x"F05A", x"F6D6",
		x"FF80", x"087C", x"0F69", x"12BF", x"1224", x"0E26", x"0805", x"0126",
		x"FA87", x"F535", x"F16C", x"EF3F", x"EE1B", x"EDB3", x"EE16", x"EF8E",
		x"F275", x"F6CF", x"FC6B", x"02D1", x"094E", x"0EF1", x"12C6", x"1440",
		x"1305", x"0F6F", x"0A47", x"042E", x"FDEB", x"F855", x"F3C9", x"F09D",
		x"EEB8", x"EDF2", x"EE05", x"EF6C", x"F23F", x"F6AA", x"FCAD", x"0387",
		x"0A65", x"0FC8", x"130C", x"137F", x"1177", x"0DCC", x"0952", x"0527",
		x"01EB", x"001C", x"FF8A", x"0041", x"0269", x"0597", x"09E8", x"0E5D",
		x"11C7", x"132B", x"11AC", x"0D28", x"062A", x"FDDB", x"F5B5", x"EF55",
		x"EC05", x"EBD4", x"EE8B", x"F300", x"F826", x"FD24", x"0146", x"0483",
		x"06CD", x"0897", x"0A74", x"0C99", x"0EEC", x"1153", x"1346", x"13E0",
		x"1252", x"0E17", x"0760", x"FF7F", x"F7D2", x"F1B4", x"EDAB", x"EBC6",
		x"EB3C", x"EB2D", x"EB10", x"EAE8", x"EABA", x"EB20", x"ED53", x"F260",
		x"FA1A", x"02E0", x"0ADD", x"1082", x"139E", x"1513", x"1573", x"1518",
		x"138D", x"101A", x"0A56", x"02CD", x"FAAB", x"F38C", x"EEF1", x"ED75",
		x"EF26", x"F3D4", x"FAC5", x"02DD", x"0AB3", x"1085", x"12DD", x"1153",
		x"0CAA", x"0632", x"FF34", x"F879", x"F299", x"EE28", x"EBFC", x"ECC8",
		x"F081", x"F6BD", x"FE80", x"066E", x"0D37", x"11DC", x"141F", x"147A",
		x"1369", x"1158", x"0E97", x"0BC7", x"0922", x"070A", x"05E2", x"055F",
		x"058F", x"0640", x"074C", x"08E8", x"0AD1", x"0D1F", x"0F5D", x"11B4",
		x"13A4", x"147F", x"13A7", x"1062", x"0AE3", x"03B4", x"FBDA", x"F4A7",
		x"EF4A", x"EC77", x"EC9D", x"EF55", x"F45C", x"FB0A", x"0260", x"096D",
		x"0F44", x"12E9", x"137E", x"106A", x"0A1F", x"0232", x"FA68", x"F3F9",
		x"EF73", x"ED15", x"EC4A", x"ECCD", x"EE75", x"F14A", x"F4E3", x"F865",
		x"FA95", x"FA5E", x"F7D4", x"F3A0", x"EFA1", x"EDBD", x"EF64", x"F466",
		x"FAC4", x"FFCD", x"0117", x"FE3A", x"F851", x"F226", x"EDFE", x"ED54",
		x"EFEB", x"F3C9", x"F67A", x"F67B", x"F3CB", x"EFE2", x"ED20", x"ED63",
		x"F132", x"F79B", x"FED7", x"0561", x"0AA5", x"0E5B", x"10CE", x"123E",
		x"12DD", x"1320", x"134D", x"1378", x"1373", x"12F6", x"11E0", x"106A",
		x"0E8D", x"0C47", x"0995", x"064F", x"028F", x"FEC6", x"FB61", x"F887",
		x"F62C", x"F460", x"F320", x"F26B", x"F249", x"F286", x"F354", x"F497",
		x"F66D", x"F8E7", x"FC85", x"0186", x"0780", x"0D5C", x"11C2", x"1376",
		x"11E7", x"0D7B", x"0765", x"015B", x"FD1A", x"FB4A", x"FBF7", x"FEA4",
		x"028D", x"06BD", x"0A6E", x"0CF3", x"0D70", x"0B91", x"070B", x"007E",
		x"F90B", x"F234", x"EDB2", x"EC49", x"EDBE", x"F117", x"F4BD", x"F7DD",
		x"F9B5", x"FAE6", x"FC36", x"FE51", x"019C", x"060A", x"0B0A", x"0FA1",
		x"12A1", x"12B7", x"0FAD", x"0A2E", x"03F6", x"FEBD", x"FB58", x"FA31",
		x"FB24", x"FDA5", x"010F", x"04D6", x"086C", x"0B8C", x"0E26", x"1028",
		x"11C6", x"12DC", x"13AE", x"1430", x"149D", x"14B9", x"1409", x"11F0",
		x"0DEC", x"07FB", x"00AF", x"F92C", x"F28F", x"EDD2", x"EBD7", x"ED1C",
		x"F16F", x"F825", x"FFFD", x"07A6", x"0DE0", x"121C", x"1427", x"1478",
		x"13C4", x"12A8", x"11BF", x"10F6", x"1003", x"0E8E", x"0BF7", x"07D7",
		x"01DA", x"FAA5", x"F38F", x"EE8E", x"ECE1", x"EE4F", x"F12B", x"F36C",
		x"F381", x"F18F", x"EED2", x"EDBD", x"EFE3", x"F56F", x"FC7B", x"0248",
		x"046B", x"01E0", x"FBB6", x"F461", x"EED8", x"ED39", x"EF0A", x"F241",
		x"F41E", x"F35E", x"F0BC", x"EE22", x"EDF4", x"F129", x"F756", x"FE2C",
		x"0318", x"043F", x"015B", x"FBB1", x"F53C", x"EFD4", x"ED16", x"EDDC",
		x"F1AC", x"F73C", x"FCD8", x"016D", x"049C", x"06C2", x"0855", x"0993",
		x"0A5A", x"0AAB", x"0A5C", x"0950", x"078C", x"0503", x"01F9", x"FECF",
		x"FBBC", x"F8B5", x"F5C0", x"F301", x"F0BE", x"EF08", x"EDC2", x"ECAD",
		x"EBAA", x"EB06", x"EABF", x"EAB2", x"EAD4", x"EB1D", x"EB7D", x"EC3F",
		x"ED83", x"F004", x"F408", x"F9F0", x"0135", x"08DD", x"0F21", x"127D",
		x"12F8", x"115A", x"0F15", x"0D9F", x"0D64", x"0E91", x"1075", x"12B3",
		x"144E", x"1543", x"15A3", x"156E", x"141C", x"1138", x"0C77", x"05A8",
		x"FD9C", x"F580", x"EF2B", x"EC0E", x"EC62", x"EFB6", x"F522", x"FBDB",
		x"0322", x"0A0C", x"0FC6", x"1305", x"1351", x"1084", x"0ADD", x"034B",
		x"FB41", x"F43D", x"EF38", x"EC5C", x"EAFE", x"EA91", x"EA89", x"EB05",
		x"EC05", x"EDE2", x"F04F", x"F328", x"F608", x"F89B", x"FAB4", x"FC21",
		x"FD22", x"FE43", x"0063", x"03DF", x"0899", x"0DA0", x"1180", x"12F1",
		x"10E5", x"0BC3", x"0524", x"FED8", x"FAAB", x"F9A9", x"FC0F", x"0108",
		x"0767", x"0D6B", x"119A", x"130F", x"1154", x"0D2C", x"0796", x"01DF",
		x"FCD6", x"F8C6", x"F5FB", x"F489", x"F4AC", x"F692", x"FA6D", x"0045",
		x"0761", x"0E08", x"1254", x"1351", x"11E0", x"0FB1", x"0EC9", x"0FB5",
		x"119D", x"12B8", x"1106", x"0BFA", x"045F", x"FCBB", x"F727", x"F4DE",
		x"F5D6", x"F933", x"FDF4", x"02B1", x"06A5", x"08FC", x"08F6", x"05FC",
		x"0064", x"F940", x"F27D", x"EE02", x"ECB5", x"EE14", x"F0C9", x"F378",
		x"F507", x"F4E3", x"F34A", x"F0FA", x"EE8A", x"EC5D", x"EADC", x"EA2D",
		x"EA60", x"EB3F", x"ECA9", x"EE47", x"F005", x"F1A3", x"F2C1", x"F32F",
		x"F2D6", x"F1F1", x"F08B", x"EED9", x"ED43", x"EBF2", x"EB20", x"EAA3",
		x"EA78", x"EAA6", x"EAEA", x"EB76", x"EC34", x"ED82", x"EF59", x"F19E",
		x"F3F8", x"F647", x"F849", x"F9EF", x"FB84", x"FD3A", x"FF7B", x"02AF",
		x"06F1", x"0BF3", x"1059", x"12F3", x"12A1", x"0F45", x"09CC", x"035A",
		x"FD71", x"F942", x"F75B", x"F7A7", x"F9AE", x"FCF1", x"00DB", x"04F6",
		x"08C0", x"0BC8", x"0E2A", x"0FCD", x"10D1", x"11BA", x"12BF", x"13E6",
		x"14D2", x"1502", x"13D2", x"10E5", x"0C21", x"05B1", x"FE60", x"F71C",
		x"F103", x"ED2A", x"EC9B", x"EFBE", x"F5F4", x"FDDA", x"05D3", x"0CA4",
		x"1182", x"1458", x"157C", x"159F", x"1577", x"1573", x"1585", x"1538",
		x"1433", x"11FA", x"0E2A", x"0839", x"005F", x"F7F5", x"F0DF", x"ECCD",
		x"EBFB", x"ED5A", x"EF0B", x"EF70", x"EE4F", x"ED05", x"ED58", x"F0C1",
		x"F6FE", x"FEE6", x"0603", x"0A18", x"098E", x"049E", x"FCE9", x"F503",
		x"EF32", x"ECE0", x"ED6D", x"EF87", x"F160", x"F1D0", x"F0BA", x"EEC9",
		x"ED0F", x"EBB2", x"EAE7", x"EA68", x"EA6F", x"EB92", x"EE69", x"F358",
		x"FA3B", x"0264", x"0A3D", x"1041", x"13A7", x"14D5", x"1492", x"136A",
		x"121B", x"10E3", x"1035", x"0FD1", x"0FA7", x"0F7A", x"0FAB", x"1063",
		x"1189", x"12A9", x"13B2", x"145E", x"14A6", x"146B", x"1398", x"1247",
		x"1083", x"0EC9", x"0CF4", x"0B8A", x"0A4A", x"094F", x"0906", x"0931",
		x"09FD", x"0B4A", x"0D3D", x"0F9B", x"1203", x"13FE", x"147F", x"12FD",
		x"0F24", x"08F6", x"01A9", x"FA54", x"F3DF", x"EEF9", x"EBFA", x"EAEC",
		x"EB96", x"ED4B", x"EF6A", x"F12B", x"F1EA", x"F159", x"EFB7", x"EDAB",
		x"EC40", x"EC77", x"EF00", x"F425", x"FB5C", x"032B", x"0A06", x"0F06",
		x"1209", x"138C", x"1425", x"1456", x"1478", x"14A1", x"1465", x"1322",
		x"0F8F", x"0942", x"00D6", x"F835", x"F134", x"ECCB", x"EAAC", x"E9FD",
		x"EA41", x"EBD4", x"EF41", x"F4E9", x"FCC6", x"056B", x"0D28", x"127A",
		x"1513", x"158F", x"1531", x"1478", x"13BC", x"12BE", x"115F", x"0F67",
		x"0C65", x"07E9", x"01F4", x"FAF2", x"F41F", x"EEB6", x"EC0E", x"EC9F",
		x"F071", x"F6BC", x"FE94", x"067F", x"0D3F", x"1202", x"1451", x"1435",
		x"1216", x"0E86", x"0A03", x"0526", x"007B", x"FC7C", x"F9E5", x"F92C",
		x"FAD7", x"FEB9", x"0458", x"0ABE", x"1030", x"1322", x"12D9", x"1023",
		x"0CAF", x"0A7D", x"0A50", x"0C81", x"0FD4", x"12A7", x"1321", x"1018",
		x"09B3", x"00F0", x"F7EB", x"F0C1", x"ECFA", x"ED28", x"F0AB", x"F616",
		x"FB76", x"FF11", x"FFA2", x"FCED", x"F7D5", x"F21E", x"EDE1", x"ECBD",
		x"EEDE", x"F323", x"F7AE", x"FB20", x"FC3C", x"FB28", x"F866", x"F4DD",
		x"F161", x"EE98", x"EC83", x"EB45", x"EAD1", x"EAEF", x"EBBC", x"ECDB",
		x"EE11", x"EEB3", x"EEAE", x"EDCF", x"ECCA", x"EC60", x"EDB5", x"F17A",
		x"F7C1", x"FFB4", x"0793", x"0DC4", x"11CC", x"1415", x"1527", x"1577",
		x"158F", x"157D", x"1536", x"147F", x"1346", x"1169", x"0EBE", x"0BA5",
		x"084C", x"0583", x"0414", x"0471", x"0713", x"0B33", x"0FB5", x"12F5",
		x"1334", x"1010", x"0A6F", x"0458", x"FFD2", x"FDE3", x"FEB5", x"019D",
		x"05A5", x"09B9", x"0CF0", x"0ED6", x"0F0C", x"0D7F", x"0A28", x"04D2",
		x"FDEC", x"F689", x"F04C", x"ECCE", x"ED2D", x"F17A", x"F8AC", x"010B",
		x"08F4", x"0F0D", x"12B2", x"1409", x"13B8", x"12D0", x"1202", x"1202",
		x"12C1", x"13DB", x"14BA", x"14FC", x"14BB", x"1437", x"13E7", x"13F5",
		x"1455", x"14A5", x"14B4", x"143C", x"1360", x"120D", x"1097", x"0EFC",
		x"0D79", x"0C3D", x"0AF4", x"094B", x"06A0", x"0290", x"FD36", x"F769",
		x"F1D1", x"EDF0", x"EC9A", x"EE71", x"F2CF", x"F826", x"FCCB", x"FF88",
		x"000D", x"FE92", x"FBBA", x"F82C", x"F49A", x"F172", x"EF45", x"EE87",
		x"EF63", x"F1AB", x"F4FC", x"F8BE", x"FC3B", x"FEB3", x"FF8C", x"FE77",
		x"FB81", x"F709", x"F22E", x"EE1D", x"EC42", x"ED79", x"F242", x"F9DE",
		x"02CF", x"0B4D", x"1169", x"1415", x"1351", x"1016", x"0BBA", x"077E",
		x"048F", x"02FD", x"02E1", x"0422", x"0691", x"09C6", x"0D32", x"102A",
		x"126C", x"1408", x"14EF", x"1557", x"1535", x"14BA", x"13FF", x"133D",
		x"12D5", x"12E0", x"136E", x"142E", x"14B3", x"14A1", x"13FD", x"1352",
		x"132E", x"13A1", x"13FE", x"130E", x"0FCB", x"09EC", x"0215", x"F9F8",
		x"F350", x"EF52", x"EDF0", x"EE9F", x"F0F0", x"F440", x"F823", x"FBC9",
		x"FE0E", x"FE17", x"FBA0", x"F726", x"F1ED", x"EE1A", x"ED1F", x"EF5D",
		x"F3E8", x"F909", x"FD2A", x"FF27", x"FF03", x"FD1E", x"FA29", x"F6D5",
		x"F376", x"F06E", x"EDD7", x"EC17", x"EB0F", x"EABC", x"EAF6", x"EB54",
		x"EBD3", x"EC37", x"EC78", x"EC85", x"EC4B", x"EBF3", x"EB94", x"EB5E",
		x"EB6B", x"EBD9", x"ECA4", x"EDD8", x"EF6C", x"F12F", x"F32A", x"F557",
		x"F79C", x"F9FB", x"FC4D", x"FEAC", x"0106", x"0363", x"05A0", x"07AA",
		x"0962", x"0B3E", x"0DCC", x"10B7", x"1329", x"13E0", x"1209", x"0D61",
		x"06B0", x"FF27", x"F81A", x"F2CC", x"EFAB", x"EE81", x"EE75", x"EF48",
		x"F110", x"F3E3", x"F80C", x"FD0F", x"0287", x"0818", x"0D40", x"1176",
		x"13BF", x"1377", x"1024", x"0A3F", x"02BE", x"FAE1", x"F3EF", x"EEEC",
		x"EC43", x"EBFB", x"EE4E", x"F319", x"FA14", x"0217", x"09AE", x"0F85",
		x"1287", x"12A3", x"100F", x"0BAF", x"06C0", x"028C", x"FFBA", x"FE79",
		x"FEC4", x"009D", x"03CD", x"07E8", x"0C70", x"1067", x"1336", x"144F",
		x"137C", x"1086", x"0BB6", x"056B", x"FE29", x"F6AA", x"F08E", x"EDB2",
		x"EED3", x"F3E9", x"FB1F", x"028B", x"08A7", x"0CA6", x"0DE6", x"0C6E",
		x"087F", x"0280", x"FB86", x"F491", x"EF2F", x"EC98", x"ED32", x"F074",
		x"F522", x"F9EB", x"FDD1", x"0062", x"019B", x"0173", x"0012", x"FD45",
		x"F976", x"F4E3", x"F081", x"ED65", x"EC80", x"EE95", x"F3C8", x"FB8B",
		x"0429", x"0BF9", x"115D", x"139F", x"1325", x"10AD", x"0D2D", x"0988",
		x"0696", x"04AF", x"0409", x"04BE", x"06CB", x"0A01", x"0DA9", x"1115",
		x"134A", x"138C", x"1128", x"0C05", x"04E2", x"FD2C", x"F678", x"F196",
		x"EE72", x"ECC4", x"EC0B", x"EC0D", x"ECC0", x"EE3F", x"F11C", x"F553",
		x"FAD3", x"0161", x"084A", x"0E87", x"127F", x"1369", x"116E", x"0DA9",
		x"09D2", x"0716", x"060D", x"0707", x"098C", x"0CA8", x"0FB9", x"1227",
		x"13A3", x"13C0", x"11D4", x"0D9B", x"070F", x"FF3C", x"F72C", x"F07D",
		x"EC76", x"EB65", x"EC85", x"EE70", x"F024", x"F166", x"F254", x"F3A1",
		x"F5B3", x"F90E", x"FDF8", x"0430", x"0AC0", x"104E", x"1390", x"13EB",
		x"1171", x"0CCC", x"075C", x"0222", x"FDD7", x"FA7F", x"F7DF", x"F595",
		x"F3CF", x"F26F", x"F156", x"F033", x"EEF4", x"EDC1", x"ECAB", x"EBFF",
		x"EB6B", x"EB13", x"EB6D", x"ECE5", x"F01B", x"F511", x"FB88", x"02DA",
		x"0A0B", x"0FF5", x"135C", x"137B", x"108A", x"0B3D", x"0495", x"FD38",
		x"F62F", x"F081", x"ED13", x"EC2E", x"EE17", x"F24D", x"F896", x"FFE6",
		x"070C", x"0D41", x"11DB", x"1420", x"1300", x"0E59", x"06B5", x"FDDE",
		x"F5AA", x"EFAA", x"EC06", x"EA4F", x"E9F3", x"EADD", x"ED81", x"F24E",
		x"F916", x"010C", x"0908", x"0FAB", x"1380", x"13E2", x"1093", x"0A58",
		x"0247", x"F9E9", x"F29C", x"ED8C", x"EAD7", x"EA1D", x"EA9E", x"EC2A",
		x"EF42", x"F4D0", x"FCC1", x"0599", x"0D74", x"122E", x"1345", x"10DF",
		x"0BF2", x"057D", x"FE13", x"F6F7", x"F138", x"ED7A", x"EB9D", x"EB09",
		x"EB60", x"EC13", x"ED2B", x"EE26", x"EF31", x"F05B", x"F1B1", x"F36D",
		x"F599", x"F862", x"FB94", x"FEE4", x"0227", x"0508", x"0759", x"0908",
		x"0A56", x"0B8C", x"0CE3", x"0E8E", x"107C", x"1285", x"1413", x"1462",
		x"1308", x"0FC2", x"0AB6", x"042A", x"FCCA", x"F585", x"EFB2", x"ECB5",
		x"EDD7", x"F2EE", x"FAF4", x"0392", x"0B20", x"1086", x"13A4", x"1495",
		x"12D5", x"0E69", x"076B", x"FF27", x"F725", x"F0CC", x"ECBF", x"EAA0",
		x"EA48", x"EB05", x"ED25", x"F120", x"F776", x"FFDE", x"08B7", x"0FDE",
		x"1345", x"11F0", x"0C8D", x"0499", x"FC3B", x"F518", x"F00C", x"ED21",
		x"EC22", x"ED2F", x"F056", x"F5B6", x"FCC8", x"04B1", x"0C13", x"11B5",
		x"14C1", x"1575", x"1517", x"14D5", x"14D3", x"1476", x"1314", x"10AC",
		x"0DCE", x"0B35", x"0914", x"076D", x"062E", x"04DA", x"0303", x"0012",
		x"FC38", x"F7AD", x"F301", x"EF19", x"ECFE", x"ED91", x"F0F1", x"F67B",
		x"FCFF", x"036C", x"0901", x"0D20", x"0FF7", x"1195", x"1289", x"1341",
		x"13E3", x"1462", x"14C5", x"14D1", x"142D", x"12D1", x"10CD", x"0E8D",
		x"0CD8", x"0C77", x"0DE0", x"1035", x"1218", x"1203", x"0F0A", x"0960",
		x"0232", x"FB8B", x"F779", x"F786", x"FBDF", x"02FB", x"0A8E", x"1041",
		x"12E6", x"12E0", x"1165", x"103C", x"1087", x"121E", x"139F", x"12F3",
		x"0EDD", x"07CF", x"FEF2", x"F649", x"EFC6", x"EC90", x"ED17", x"F0E7",
		x"F6D3", x"FD31", x"031A", x"07A2", x"0A2E", x"0A91", x"08E4", x"05B5",
		x"01CD", x"FDCF", x"FA5A", x"F7FE", x"F6F8", x"F787", x"F980", x"FC7B",
		x"FFCB", x"0310", x"0604", x"0868", x"09FE", x"0A72", x"09F0", x"0893",
		x"0696", x"03D7", x"0042", x"FBE2", x"F737", x"F29F", x"EEBA", x"EC7E",
		x"ECA6", x"EF9A", x"F4DA", x"FB6F", x"023C", x"0865", x"0D6E", x"10F9",
		x"1346", x"1488", x"152F", x"1559", x"1524", x"14CF", x"1476", x"142C",
		x"13A0", x"128B", x"10F3", x"0F31", x"0D95", x"0C5D", x"0BC6", x"0BCA",
		x"0C2F", x"0D01", x"0E49", x"102E", x"1267", x"1409", x"13EE", x"113A",
		x"0BBC", x"0411", x"FBD2", x"F47B", x"EEFD", x"EBB9", x"EA87", x"EB25",
		x"ED6C", x"F1AB", x"F7EC", x"FFFC", x"0873", x"0F78", x"139E", x"14CD",
		x"13E5", x"1219", x"1042", x"0EEE", x"0E29", x"0DD2", x"0DB9", x"0DAD",
		x"0DB6", x"0DE2", x"0E5E", x"0F6A", x"10F6", x"12BA", x"13F2", x"1412",
		x"1249", x"0E1E", x"07A7", x"FFBE", x"F7EA", x"F19E", x"ED5D", x"EB3C",
		x"EA9F", x"EAC5", x"EB66", x"EC8D", x"EE5F", x"F0B3", x"F2B3", x"F344",
		x"F24F", x"F025", x"EE04", x"ED9B", x"F012", x"F5B9", x"FD21", x"0411",
		x"08AE", x"0A41", x"0959", x"0696", x"02B1", x"FE17", x"FA09", x"F798",
		x"F7A4", x"FA8D", x"FFF4", x"06E1", x"0D6B", x"11DD", x"133C", x"11D7",
		x"0EF8", x"0BFB", x"0A10", x"09C2", x"0B25", x"0DBE", x"1077", x"12AA",
		x"141F", x"14E7", x"1516", x"14F4", x"146D", x"1397", x"1270", x"10F8",
		x"0F46", x"0D30", x"0ADD", x"085F", x"05CA", x"0343", x"00D1", x"FE63",
		x"FC21", x"F9FC", x"F7C7", x"F54C", x"F2D2", x"F0C6", x"EF04", x"ED89",
		x"EC46", x"EB54", x"EAF7", x"EB15", x"EB48", x"EB76", x"EB93", x"EBF4",
		x"ECD2", x"EEAA", x"F218", x"F772", x"FEA1", x"06BC", x"0E08", x"12D4",
		x"146C", x"1381", x"11A3", x"109B", x"1115", x"1283", x"1367", x"120D",
		x"0D91", x"064C", x"FD80", x"F539", x"EF27", x"EC09", x"EC0A", x"EED1",
		x"F3AF", x"FA50", x"01A7", x"08CA", x"0E99", x"1253", x"1375", x"120A",
		x"0E99", x"093E", x"026E", x"FADD", x"F3D3", x"EECD", x"ED0D", x"EECA",
		x"F378", x"FA12", x"00F9", x"06A7", x"0A1E", x"0B2E", x"0A4D", x"07D4",
		x"047F", x"00D8", x"FDA2", x"FB5B", x"FAD2", x"FC5C", x"003C", x"05B9",
		x"0B9F", x"1047", x"1241", x"111C", x"0CB2", x"05F1", x"FE34", x"F6C0",
		x"F0EB", x"ED44", x"EC11", x"ED49", x"F130", x"F74B", x"FF08", x"070F",
		x"0E05", x"1292", x"1432", x"132C", x"1015", x"0BAC", x"069E", x"017C",
		x"FCE5", x"F93D", x"F699", x"F4F1", x"F41C", x"F3E4", x"F3EF", x"F446",
		x"F4E0", x"F5C9", x"F728", x"F912", x"FC19", x"008B", x"063F", x"0C13",
		x"10A5", x"12BE", x"119E", x"0DBD", x"082A", x"02D3", x"FF41", x"FEA4",
		x"0122", x"05E2", x"0B94", x"1058", x"12B1", x"1182", x"0CB3", x"04F7",
		x"FBF2", x"F3B2", x"EE23", x"EBFC", x"ECFB", x"F01F", x"F400", x"F731",
		x"F897", x"F800", x"F5CC", x"F2F7", x"F051", x"EE33", x"ECB1", x"EC00",
		x"ED0C", x"F09A", x"F6DD", x"FECB", x"06E8", x"0DC1", x"127A", x"14E1",
		x"156E", x"153F", x"14EF", x"14A9", x"13F3", x"12A6", x"112B", x"106A",
		x"10DF", x"1207", x"1349", x"131D", x"10C5", x"0B9D", x"0489", x"FCA2",
		x"F5AF", x"F075", x"ED0E", x"EB6E", x"EAF5", x"EAED", x"EAE5", x"EAF1",
		x"EB07", x"EB3C", x"EB39", x"EB2E", x"EAF7", x"EB05", x"EB9B", x"ECA1",
		x"EE22", x"EFFB", x"F21D", x"F45C", x"F6D2", x"F97C", x"FC27", x"FF03",
		x"018C", x"03BF", x"0591", x"0716", x"08B1", x"0A58", x"0C1E", x"0E32",
		x"1076", x"12B2", x"1442", x"146B", x"1261", x"0DFD", x"0782", x"FFFE",
		x"F8AB", x"F2AC", x"EE69", x"EBFD", x"EB56", x"EBF0", x"ED1F", x"EE5B",
		x"EF18", x"EEFE", x"EE17", x"ECDA", x"EBD0", x"EBE5", x"EDF3", x"F268",
		x"F973", x"01C8", x"09DA", x"1002", x"138A", x"1420", x"1213", x"0DE7",
		x"07E3", x"00E2", x"F98C", x"F2DD", x"EE60", x"ED4C", x"F01E", x"F61C",
		x"FD95", x"04C3", x"0A5C", x"0D4B", x"0D14", x"09A6", x"03B9", x"FC6A",
		x"F554", x"EFCE", x"ECF9", x"ED2B", x"EF68", x"F27C", x"F526", x"F709",
		x"F80A", x"F8F9", x"FA9E", x"FDD5", x"02B8", x"0885", x"0E0E", x"11D8",
		x"12CE", x"1097", x"0BE6", x"069A", x"02E7", x"026C", x"0573", x"0AA4",
		x"0FDF", x"12ED", x"1276", x"0E9A", x"08B9", x"0263", x"FD18", x"F9B6",
		x"F7F1", x"F740", x"F67E", x"F4ED", x"F256", x"EF60", x"ED1C", x"ED1F",
		x"F046", x"F631", x"FDCA", x"053B", x"0B04", x"0E19", x"0E22", x"0AE4",
		x"0508", x"FDBF", x"F674", x"F08C", x"ED07", x"EC7F", x"EE8F", x"F258",
		x"F6F9", x"FB72", x"FF20", x"01CE", x"02EC", x"0212", x"FF3D", x"FA80",
		x"F4BC", x"EFBF", x"ED1B", x"EDD8", x"F13F", x"F5C4", x"F907", x"F9CB",
		x"F7B1", x"F385", x"EF38", x"ECFF", x"EE0A", x"F271", x"F902", x"0033",
		x"069B", x"0BA3", x"0F1D", x"1156", x"12B4", x"1337", x"12D9", x"1139",
		x"0DE4", x"0885", x"0197", x"FA0B", x"F34B", x"EE89", x"EC00", x"EB62",
		x"EBCE", x"EC8C", x"EC9F", x"EC15", x"EB62", x"EB04", x"EB4F", x"EC93",
		x"EE89", x"F0FC", x"F3F6", x"F75B", x"FACD", x"FDC2", x"FF7D", x"FF54",
		x"FD42", x"F96A", x"F4A2", x"EFDC", x"ED03", x"ED05", x"F01D", x"F50E",
		x"FA30", x"FE0D", x"FFD3", x"FF3B", x"FCD1", x"F949", x"F552", x"F18B",
		x"EE71", x"EC9F", x"EBBC", x"EB7A", x"EB28", x"EADD", x"EABA", x"EB0B",
		x"EC17", x"EE6A", x"F2AA", x"F90F", x"00EE", x"08EE", x"0F79", x"1372",
		x"14DD", x"1499", x"13E2", x"1396", x"13D1", x"144A", x"148E", x"14C3",
		x"1483", x"13E5", x"1347", x"12FE", x"1314", x"1389", x"1430", x"14AE",
		x"14D5", x"141D", x"11C5", x"0D29", x"063C", x"FDF0", x"F5E5", x"EFD8",
		x"EC6D", x"EB29", x"EAF0", x"EB11", x"EB83", x"ED3B", x"F117", x"F770",
		x"FF80", x"07A8", x"0E3F", x"120A", x"137C", x"1320", x"11DE", x"0FE6",
		x"0D2C", x"0997", x"057C", x"016E", x"FD9F", x"FA05", x"F696", x"F377",
		x"F0F4", x"EF2D", x"EE62", x"EEEA", x"F177", x"F660", x"FD7D", x"0569",
		x"0C84", x"118B", x"13F0", x"1418", x"131E", x"124C", x"1239", x"1312",
		x"1419", x"14B1", x"1488", x"1402", x"139A", x"13D1", x"146C", x"14C5",
		x"1464", x"137F", x"1285", x"120B", x"1251", x"1315", x"1377", x"125F",
		x"0EF9", x"0907", x"0168", x"F9A7", x"F373", x"EFD6", x"EEF5", x"EFF9",
		x"F256", x"F579", x"F8EE", x"FC46", x"FEF9", x"009C", x"0122", x"0079",
		x"FE92", x"FBAE", x"F886", x"F567", x"F2CD", x"F096", x"EEC4", x"ED4C",
		x"EC02", x"EB32", x"EAEC", x"EB32", x"EBBA", x"EC02", x"EBF1", x"EB86",
		x"EB26", x"EAE6", x"EB46", x"EC34", x"ED52", x"EE2E", x"EE5D", x"EE34",
		x"EDB0", x"ED18", x"EC55", x"EB8A", x"EB28", x"EB3D", x"EBE5", x"ED11",
		x"EEF2", x"F1BA", x"F4ED", x"F83C", x"FAD8", x"FC36", x"FBE8", x"F9B8",
		x"F5E7", x"F17E", x"EDEF", x"ECB2", x"EEBC", x"F364", x"F998", x"FFFB",
		x"059C", x"09F6", x"0CD1", x"0E99", x"0FFF", x"116B", x"12C6", x"13DC",
		x"1487", x"14C9", x"14E7", x"14F3", x"14DA", x"147C", x"13A9", x"11C6",
		x"0E71", x"0948", x"0276", x"FAFC", x"F412", x"EEEA", x"EC2E", x"EC0B",
		x"EE2C", x"F208", x"F6D1", x"FB8A", x"FF8F", x"0247", x"0374", x"0338",
		x"017B", x"FE6F", x"FA12", x"F50B", x"F056", x"ED1D", x"EC6B", x"EEEF",
		x"F4C3", x"FCE3", x"05DD", x"0D7B", x"1245", x"1376", x"1143", x"0D6E",
		x"0A24", x"08F2", x"0A6B", x"0DDD", x"1165", x"12E9", x"10FB", x"0C0A",
		x"05E8", x"012A", x"FFBC", x"0216", x"0743", x"0CF3", x"1101", x"11E9",
		x"0F7B", x"0A92", x"04C0", x"FF81", x"FBFD", x"FA55", x"F9B8", x"F92C",
		x"F79A", x"F4C4", x"F12B", x"EE1F", x"ECC0", x"EDDC", x"F1E1", x"F7E6",
		x"FEFC", x"05AE", x"0ACE", x"0DE4", x"0ED1", x"0E20", x"0C1D", x"091E",
		x"0581", x"017C", x"FD74", x"F9DF", x"F74C", x"F58D", x"F45A", x"F342",
		x"F201", x"F04E", x"EE51", x"EC86", x"EC43", x"EEAE", x"F418", x"FBA7",
		x"03AD", x"0AAD", x"0FD7", x"1291", x"12B1", x"105F", x"0BC1", x"0518",
		x"FD08", x"F517", x"EEBC", x"EB9C", x"EB89", x"ED7F", x"EFAF", x"F107",
		x"F1A5", x"F227", x"F349", x"F5A7", x"F9E1", x"000B", x"0777", x"0E55",
		x"12B1", x"135D", x"10F2", x"0D89", x"0B06", x"0AEE", x"0D28", x"1089",
		x"12D6", x"1226", x"0DF4", x"076A", x"00C2", x"FC18", x"FA7B", x"FBE3",
		x"FFA5", x"0475", x"08D3", x"0C11", x"0DB3", x"0D3E", x"09B1", x"0304",
		x"FAA7", x"F316", x"EE41", x"ECAB", x"ED2C", x"EE03", x"EE27", x"ED68",
		x"ECC3", x"ED90", x"F0FD", x"F720", x"FF0B", x"06DC", x"0D40", x"11B0",
		x"142B", x"1545", x"1575", x"156E", x"154F", x"1553", x"1566", x"1561",
		x"1542", x"14F5", x"141B", x"12E1", x"1189", x"1067", x"0FAD", x"0F81",
		x"0FE3", x"10AA", x"11BC", x"12D3", x"13B7", x"1450", x"148E", x"1444",
		x"134C", x"1185", x"0EEC", x"0BE8", x"0945", x"07CF", x"07D1", x"0995",
		x"0CC1", x"102C", x"12A6", x"12D8", x"0FD2", x"0A2D", x"0374", x"FDAA",
		x"FA2E", x"F956", x"FABE", x"FDB8", x"018C", x"0551", x"0851", x"0A9B",
		x"0BFB", x"0C6B", x"0BE8", x"0A5C", x"081D", x"0533", x"0177", x"FCE3",
		x"F7DC", x"F2ED", x"EECE", x"EC62", x"EC81", x"EF5B", x"F4A1", x"FB36",
		x"0205", x"07FB", x"0CB6", x"101C", x"1262", x"13B7", x"1482", x"14EF",
		x"1502", x"14EB", x"14A6", x"13FC", x"12F3", x"11AD", x"1035", x"0E60",
		x"0BFE", x"08F1", x"056D", x"0182", x"FD6D", x"F96C", x"F5EF", x"F3A7",
		x"F326", x"F4A0", x"F86E", x"FE5B", x"058D", x"0C6E", x"1114", x"12F4",
		x"1269", x"10EF", x"1056", x"110E", x"128C", x"135A", x"11F0", x"0D75",
		x"067D", x"FE88", x"F72D", x"F140", x"ED6A", x"EB73", x"EAFC", x"EB2E",
		x"EB52", x"EB1D", x"EADE", x"EB3F", x"ED31", x"F11F", x"F729", x"FE92",
		x"064F", x"0D0E", x"11F1", x"1490", x"14E7", x"13ED", x"1232", x"1037",
		x"0E60", x"0CFC", x"0C72", x"0CFE", x"0E8B", x"107D", x"1269", x"13F4",
		x"14CE", x"1514", x"1506", x"14EE", x"1450", x"1246", x"0E40", x"07F9",
		x"005F", x"F8A8", x"F20D", x"ED99", x"EB6B", x"EAD9", x"EAEB", x"EAEF",
		x"EB43", x"EC78", x"EEF6", x"F2CF", x"F7BA", x"FDC6", x"049D", x"0B41",
		x"107A", x"1366", x"13A0", x"117B", x"0D9F", x"08A6", x"03AC", x"FF3F",
		x"FBB6", x"F926", x"F768", x"F676", x"F655", x"F6EE", x"F819", x"F9D3",
		x"FC00", x"FEA4", x"017C", x"045A", x"06A1", x"0868", x"0968", x"094E",
		x"082E", x"05B0", x"0258", x"FE3A", x"F9EF", x"F57B", x"F158", x"EE06",
		x"EC25", x"EC5F", x"EF25", x"F462", x"FB77", x"037B", x"0B03", x"10A6",
		x"138D", x"1376", x"1091", x"0B8B", x"0552", x"FEC3", x"F894", x"F39A",
		x"EFF6", x"ED95", x"EC2C", x"EB69", x"EB08", x"EB16", x"EB29", x"EB48",
		x"EB60", x"EB6F", x"EBAF", x"EC1E", x"ED2B", x"EF20", x"F280", x"F7A5",
		x"FEA4", x"06A6", x"0DD2", x"124D", x"1359", x"11D2", x"0F7D", x"0E3C",
		x"0EE6", x"10F1", x"128C", x"11C8", x"0D7E", x"0690", x"FF66", x"FA63",
		x"F979", x"FD09", x"03B5", x"0AFD", x"1086", x"12D5", x"11D2", x"0EFC",
		x"0C33", x"0AE2", x"0BC1", x"0E2E", x"1105", x"1359", x"14D9", x"15BF",
		x"15AF", x"140B", x"0FFB", x"09A1", x"01D2", x"F9D0", x"F305", x"EE07",
		x"EB40", x"EA4C", x"EA76", x"EB10", x"EBD7", x"ED08", x"EEC1", x"F0B6",
		x"F277", x"F35C", x"F355", x"F269", x"F0CF", x"EF2C", x"ED78", x"EC38",
		x"EB78", x"EB1D", x"EB58", x"EC09", x"ED45", x"EEF8", x"F0FC", x"F2E3",
		x"F451", x"F513", x"F53B", x"F49F", x"F373", x"F1B4", x"EFA4", x"EDB3",
		x"EC2F", x"EB48", x"EAFD", x"EB23", x"EB59", x"EBC0", x"EC68", x"ED59",
		x"EE95", x"F052", x"F294", x"F57D", x"F913", x"FD25", x"0126", x"049B",
		x"0712", x"07F1", x"06DC", x"0397", x"FE4E", x"F7E2", x"F1F3", x"EE00",
		x"ECFB", x"EEC9", x"F2AA", x"F744", x"FBC5", x"FF85", x"0222", x"03E1",
		x"0576", x"0776", x"0A1E", x"0D44", x"106F", x"12B4", x"1387", x"1211",
		x"0DD5", x"0715", x"FF04", x"F718", x"F0CF", x"ED0D", x"EC2D", x"EE25",
		x"F268", x"F859", x"FEF1", x"0586", x"0B4C", x"0FE4", x"12FB", x"14B0",
		x"157D", x"15B3", x"15BC", x"1597", x"156E", x"14C1", x"132D", x"0FBD",
		x"0A3C", x"02BB", x"FA54", x"F2BE", x"EDA9", x"EC23", x"EE0A", x"F2B3",
		x"F8B8", x"FF4A", x"05D7", x"0BDE", x"10D0", x"1370", x"12A8", x"0DF6",
		x"0642", x"FD61", x"F565", x"EFC8", x"ECB8", x"EC04", x"ED92", x"F16A",
		x"F768", x"FEE8", x"06B5", x"0D68", x"1222", x"1494", x"1525", x"14C8",
		x"145F", x"1469", x"14B9", x"1495", x"1342", x"1043", x"0B3D", x"0470",
		x"FC8E", x"F4EF", x"EF30", x"EC30", x"EBE4", x"ED14", x"EE5F", x"EE84",
		x"ED8B", x"ECAE", x"EDDA", x"F237", x"F9A8", x"024B", x"09F8", x"0F64",
		x"129A", x"1441", x"1500", x"1535", x"1528", x"151B", x"14C6", x"141B",
		x"12F4", x"111C", x"0E80", x"0B62", x"088C", x"06C0", x"06C1", x"08A8",
		x"0BF7", x"0FD6", x"12E7", x"141E", x"1281", x"0E08", x"0761", x"FFEC",
		x"F913", x"F395", x"EFBE", x"ED54", x"EC0F", x"EB80", x"EB46", x"EB7F",
		x"ECF8", x"F099", x"F6BB", x"FEB3", x"06E5", x"0DB0", x"1264", x"150E",
		x"1613", x"15A7", x"13AA", x"0FB6", x"09B1", x"01FB", x"F983", x"F1F5",
		x"ED10", x"EB1E", x"EB7A", x"ED26", x"EF97", x"F295", x"F5CC", x"F870",
		x"F94A", x"F7E5", x"F4D0", x"F105", x"EDF2", x"ED02", x"EF48", x"F480",
		x"FB72", x"024C", x"07CA", x"0BA0", x"0E21", x"0FAA", x"10B7", x"1184",
		x"1247", x"1340", x"1427", x"14CE", x"14FA", x"1493", x"1398", x"1274",
		x"1188", x"1106", x"1122", x"11BE", x"12BC", x"13F0", x"14D8", x"157A",
		x"1586", x"1533", x"14C3", x"1479", x"1496", x"14B8", x"14E1", x"14A9",
		x"1412", x"1294", x"0FE1", x"0BC2", x"0651", x"0003", x"F978", x"F333",
		x"EE78", x"EC24", x"ED2D", x"F184", x"F882", x"00EA", x"0925", x"0F9F",
		x"1382", x"14BE", x"142F", x"12D9", x"11BA", x"117A", x"11EE", x"12F6",
		x"13E9", x"1491", x"14A0", x"140D", x"12F3", x"11C7", x"10B0", x"0FC1",
		x"0EC5", x"0D72", x"0B29", x"075C", x"01DC", x"FAF4", x"F418", x"EEFC",
		x"ED3C", x"EEEB", x"F2B0", x"F688", x"F85D", x"F733", x"F38E", x"EF8A",
		x"ED3E", x"EE23", x"F27E", x"F888", x"FE35", x"019E", x"020E", x"FFBB",
		x"FBBD", x"F72C", x"F30C", x"F038", x"EF30", x"F0A1", x"F4E7", x"FBCD",
		x"0439", x"0C10", x"1180", x"1415", x"1478", x"141E", x"13CC", x"136C",
		x"1212", x"0E9D", x"0882", x"008E", x"F8A3", x"F285", x"EF2A", x"EE8B",
		x"EFED", x"F285", x"F609", x"F9FE", x"FDDE", x"0090", x"0181", x"00C0",
		x"FEBE", x"FBE9", x"F892", x"F51D", x"F222", x"F039", x"EF91", x"EFEE",
		x"F0DE", x"F254", x"F445", x"F6C7", x"F9BF", x"FD18", x"0058", x"036A",
		x"0679", x"098D", x"0C81", x"0EEC", x"10DB", x"1217", x"12B5", x"1299",
		x"11A1", x"1012", x"0DF3", x"0B45", x"0858", x"05AA", x"03AB", x"02CB",
		x"033B", x"04D2", x"075D", x"0A00", x"0C95", x"0EAE", x"1085", x"11EF",
		x"12A0", x"1288", x"11CA", x"1094", x"0EF2", x"0CA2", x"0921", x"0453",
		x"FE74", x"F850", x"F2B8", x"EE97", x"ECA6", x"ED66", x"F0A2", x"F5A5",
		x"FB6F", x"00FD", x"05BB", x"0979", x"0C2A", x"0DF2", x"0F1F", x"1000",
		x"10DA", x"11C3", x"12C4", x"13B5", x"148E", x"150D", x"14F5", x"1440",
		x"1338", x"1232", x"110F", x"1002", x"0F01", x"0DCB", x"0C24", x"098B",
		x"056D", x"FFBF", x"F95D", x"F360", x"EF00", x"ED6F", x"EECE", x"F287",
		x"F6EB", x"FA17", x"FA91", x"F853", x"F455", x"F041", x"ED73", x"ED5E",
		x"F0DE", x"F7DF", x"00E1", x"09BC", x"1058", x"1371", x"1316", x"0FF2",
		x"0B8D", x"07A1", x"05A9", x"0665", x"0974", x"0D9F", x"113B", x"12D7",
		x"1167", x"0C46", x"045F", x"FB5E", x"F350", x"EDDE", x"EC10", x"EDBC",
		x"F1C5", x"F6D0", x"FB20", x"FDDC", x"FE7C", x"FD28", x"FA4D", x"F6D7",
		x"F382", x"F0D6", x"EF30", x"EF44", x"F190", x"F694", x"FDB1", x"05AA",
		x"0CC8", x"11CA", x"13F5", x"135F", x"1107", x"0E2D", x"0BD5", x"0A2D",
		x"08F6", x"076B", x"052C", x"01BC", x"FCFF", x"F74F", x"F1D1", x"EDE2",
		x"EC9A", x"EE63", x"F2CA", x"F8CA", x"FF06", x"0463", x"08CA", x"0C33",
		x"0ED7", x"10A7", x"11D4", x"1280", x"12C6", x"12C1", x"128A", x"11F1",
		x"10B2", x"0EC0", x"0BEC", x"0847", x"0400", x"FEF2", x"F97A", x"F3FF",
		x"EF52", x"EC83", x"EC78", x"EFA3", x"F566", x"FCBA", x"0465", x"0B53",
		x"10A6", x"138F", x"13F3", x"11AE", x"0D20", x"0699", x"FEDF", x"F748",
		x"F0FA", x"ED12", x"EBFC", x"ED81", x"F125", x"F5FD", x"FB58", x"00C4",
		x"060D", x"0A8E", x"0E22", x"107A", x"117E", x"1136", x"0F68", x"0B40",
		x"04A9", x"FC7C", x"F4A1", x"EF15", x"EC77", x"EBFD", x"EC53", x"EC77",
		x"EC6A", x"ED47", x"F061", x"F5FE", x"FD9A", x"052A", x"0AFB", x"0D91",
		x"0C94", x"084B", x"01CC", x"FA4F", x"F361", x"EE8E", x"ED2B", x"F01D",
		x"F6B7", x"FF3E", x"07A0", x"0E49", x"1284", x"1469", x"146D", x"1365",
		x"120C", x"1131", x"1100", x"11A8", x"12FB", x"144D", x"14F0", x"1496",
		x"1381", x"11A6", x"0FA8", x"0D85", x"0B8A", x"09E7", x"08AF", x"07C2",
		x"071B", x"06D3", x"06DC", x"0785", x"08D9", x"0ADF", x"0DB4", x"10B3",
		x"1344", x"1465", x"1390", x"1073", x"0B53", x"048E", x"FD1C", x"F62B",
		x"F0BB", x"ED4F", x"EB9F", x"EB75", x"EC92", x"EE60", x"EFF7", x"F0C0",
		x"F02B", x"EE9D", x"ECDC", x"EC07", x"ED0D", x"F06F", x"F633", x"FD41",
		x"045C", x"0A08", x"0DA8", x"0F4E", x"0F74", x"0E81", x"0C89", x"094A",
		x"049B", x"FEB2", x"F813", x"F21B", x"EE00", x"ECEB", x"EF18", x"F3B7",
		x"F957", x"FE3A", x"00DC", x"0051", x"FC9B", x"F719", x"F161", x"EDC0",
		x"ED67", x"F06E", x"F5B8", x"FBBE", x"0109", x"04D1", x"0725", x"08AB",
		x"0A08", x"0B83", x"0CF8", x"0E4E", x"0FA1", x"10FC", x"1252", x"1382",
		x"145E", x"14FA", x"1530", x"146F", x"1206", x"0D7C", x"0707", x"FF6E",
		x"F7D0", x"F163", x"ED1D", x"EB5D", x"EBD5", x"EDE7", x"F0A3", x"F399",
		x"F674", x"F8AB", x"F9C3", x"F907", x"F674", x"F2B2", x"EF28", x"ED84",
		x"EEEF", x"F3A8", x"FA2E", x"0040", x"0343", x"01F9", x"FCD0", x"F5D0",
		x"EFF7", x"ED67", x"EEA8", x"F1F4", x"F4BB", x"F50C", x"F2D7", x"EFA3",
		x"EDE2", x"EF8A", x"F491", x"FB52", x"0116", x"03A5", x"022D", x"FD34",
		x"F686", x"F097", x"ED75", x"EDE6", x"F138", x"F63D", x"FB72", x"FFBB",
		x"02DC", x"04EE", x"066C", x"07CD", x"0953", x"0B34", x"0D4F", x"0F99",
		x"11C6", x"137A", x"148B", x"152D", x"1556", x"155C", x"1590", x"159F",
		x"156E", x"1505", x"145A", x"134C", x"11A1", x"0F3C", x"0C8A", x"0A2C",
		x"0848", x"06E4", x"05B0", x"0445", x"0202", x"FE9D", x"F9FB", x"F4AC",
		x"F00C", x"ED8B", x"EE40", x"F241", x"F87F", x"FEEE", x"036C", x"04AB",
		x"020A", x"FC72", x"F5A8", x"EFFB", x"ED07", x"ED33", x"EFE1", x"F3A7",
		x"F6E1", x"F857", x"F7B8", x"F59F", x"F2BC", x"EFCC", x"ED58", x"EC05",
		x"EC5A", x"EE47", x"F20D", x"F777", x"FE14", x"0552", x"0C1E", x"1123",
		x"134C", x"11A1", x"0C93", x"0524", x"FD12", x"F5CC", x"F05C", x"ECFE",
		x"EB60", x"EAE5", x"EB22", x"EBC3", x"ED16", x"EF1B", x"F1AE", x"F3EF",
		x"F546", x"F531", x"F3C7", x"F18D", x"EF15", x"ED0F", x"EBAC", x"EADC",
		x"EA98", x"EB1F", x"ECA4", x"EFBF", x"F4BD", x"FB82", x"035D", x"0B1B",
		x"1110", x"13C1", x"127E", x"0D7D", x"0622", x"FDFD", x"F6B2", x"F119",
		x"ED68", x"EB56", x"EA8D", x"EA61", x"EAA8", x"EB59", x"ECC6", x"EECD",
		x"F109", x"F2E9", x"F3D6", x"F399", x"F22E", x"F01B", x"EDF7", x"EC35",
		x"EB1B", x"EA8B", x"EA5E", x"EA84", x"EB40", x"EC9D", x"EE9A", x"F0F6",
		x"F316", x"F42E", x"F3A2", x"F19C", x"EEE3", x"ECF0", x"ED28", x"F058",
		x"F639", x"FD5E", x"03BE", x"0808", x"09BD", x"090D", x"065A", x"0247",
		x"FDC3", x"F9DF", x"F745", x"F606", x"F61A", x"F780", x"FA1D", x"FD72",
		x"0117", x"0469", x"06F8", x"087A", x"08ED", x"0808", x"0641", x"03D9",
		x"011F", x"FE11", x"FAF6", x"F7EE", x"F4F4", x"F211", x"EF73", x"ED85",
		x"EC3D", x"EB92", x"EB44", x"EB04", x"EAEC", x"EB05", x"EB16", x"EB25",
		x"EB90", x"EC7B", x"EE1F", x"F085", x"F349", x"F620", x"F906", x"FBEF",
		x"FEEE", x"01C4", x"041B", x"05D0", x"06D1", x"076D", x"0736", x"0667",
		x"0511", x"0320", x"0090", x"FD04", x"F89C", x"F3C6", x"EF65", x"EC8D",
		x"EC06", x"EE5B", x"F34A", x"FA0C", x"013C", x"07A3", x"0C8C", x"0FB1",
		x"11AB", x"12D1", x"1395", x"1434", x"14D3", x"1514", x"1445", x"11B4",
		x"0CDA", x"0621", x"FE49", x"F6C3", x"F08F", x"EC91", x"EAFF", x"EB6F",
		x"EC9C", x"EDCD", x"EE85", x"EF4B", x"F074", x"F2B0", x"F672", x"FBF0",
		x"030B", x"0A60", x"1037", x"132C", x"12E6", x"1091", x"0DE0", x"0C84",
		x"0D6C", x"100E", x"12CB", x"13B2", x"1111", x"0B10", x"02F1", x"FA67",
		x"F2FF", x"EDD7", x"EB79", x"EC2C", x"EF8E", x"F4F6", x"FBDB", x"0333",
		x"0A30", x"0FB7", x"1311", x"13C5", x"11C8", x"0D86", x"0750", x"0005",
		x"F88B", x"F219", x"EDB2", x"EC3B", x"EDC1", x"F1C2", x"F75F", x"FDA3",
		x"03E7", x"09A9", x"0E3C", x"119D", x"13A1", x"148C", x"14E1", x"14C2",
		x"1459", x"1311", x"104E", x"0BB6", x"0540", x"FD9B", x"F5EB", x"EFCC",
		x"EC92", x"ECD1", x"F037", x"F5C5", x"FCB5", x"040F", x"0AF2", x"1030",
		x"1328", x"1372", x"1126", x"0C95", x"0669", x"FF62", x"F866", x"F261",
		x"EE1F", x"EC6E", x"EE07", x"F2BD", x"FA1F", x"0258", x"0A19", x"0FCF",
		x"134C", x"151D", x"15AB", x"1582", x"14EF", x"145E", x"1433", x"1437",
		x"13AC", x"11AF", x"0D89", x"0776", x"FFC9", x"F80C", x"F161", x"ED1C",
		x"EB9C", x"EC12", x"ECF1", x"ED3C", x"ECC0", x"EBFB", x"EC95", x"EF9D",
		x"F5A4", x"FDF9", x"06EF", x"0E5E", x"12C1", x"13B3", x"115D", x"0CD1",
		x"06F9", x"00D2", x"FA9F", x"F500", x"F07C", x"ED50", x"EB82", x"EAF7",
		x"EB34", x"EB96", x"EBD2", x"EBB0", x"EBB8", x"ECC2", x"EF67", x"F3E2",
		x"FA46", x"01DD", x"096E", x"0F78", x"1357", x"14EB", x"14A2", x"1316",
		x"1154", x"0FFF", x"0F85", x"1016", x"114B", x"12DB", x"1429", x"1456",
		x"124A", x"0D72", x"0656", x"FDED", x"F5BE", x"EF99", x"ECB5", x"EDBF",
		x"F22F", x"F89C", x"FF74", x"0582", x"0A12", x"0D19", x"0E94", x"0ED3",
		x"0E0C", x"0C78", x"09D4", x"0606", x"00E3", x"FB06", x"F536", x"F055",
		x"ED2C", x"EC52", x"EE46", x"F29D", x"F889", x"FEE2", x"047C", x"08D4",
		x"0B87", x"0D27", x"0E10", x"0F08", x"108D", x"1293", x"143C", x"144F",
		x"11B2", x"0C6A", x"051A", x"FD10", x"F58F", x"EFF9", x"ECE9", x"EC14",
		x"ECE1", x"EE94", x"F10A", x"F42A", x"F754", x"F9A4", x"FA31", x"F884",
		x"F519", x"F0DA", x"ED83", x"EC8F", x"EEF6", x"F465", x"FC0A", x"0433",
		x"0B95", x"110C", x"13EB", x"1431", x"11DA", x"0D27", x"068F", x"FEDE",
		x"F73A", x"F112", x"ED34", x"EC50", x"EE61", x"F2B5", x"F846", x"FDE9",
		x"030E", x"074D", x"0AB9", x"0D53", x"0F1F", x"1074", x"11BB", x"12DE",
		x"13B7", x"142E", x"144D", x"1466", x"14A6", x"14E0", x"1492", x"132E",
		x"1052", x"0B73", x"0453", x"FBCA", x"F3E2", x"EE40", x"EBA2", x"EB2D",
		x"EB9A", x"EBBC", x"EB95", x"EBAD", x"ED15", x"F111", x"F7C8", x"0089",
		x"095C", x"100A", x"12D2", x"114F", x"0C27", x"04F8", x"FD5F", x"F6F2",
		x"F28F", x"F122", x"F318", x"F87A", x"0025", x"0816", x"0E8C", x"127C",
		x"141B", x"143D", x"1415", x"13C9", x"12C4", x"0FD1", x"0A30", x"023A",
		x"F996", x"F28C", x"EE86", x"EDBC", x"EF6C", x"F29D", x"F67B", x"FA85",
		x"FDE2", x"FFA9", x"FF09", x"FBD6", x"F6E0", x"F169", x"ED83", x"EC99",
		x"EF1A", x"F40F", x"FA18", x"FFD1", x"047C", x"0821", x"0ACD", x"0CCE",
		x"0E5F", x"0F8E", x"1098", x"119F", x"12BA", x"13E1", x"14CE", x"1551",
		x"1544", x"14C2", x"13C2", x"12A0", x"1136", x"0F73", x"0D3A", x"0AC0",
		x"083E", x"0607", x"0449", x"02FD", x"024D", x"0256", x"0353", x"0500",
		x"0742", x"0A24", x"0D65", x"10A4", x"132D", x"146C", x"13C8", x"113B",
		x"0CC7", x"065B", x"FEA5", x"F6C9", x"F04B", x"ECCD", x"ED60", x"F202",
		x"F94A", x"011F", x"07EE", x"0CD9", x"0F49", x"0F00", x"0BE0", x"0669",
		x"FF5B", x"F7EC", x"F168", x"ED3A", x"EC26", x"EDDF", x"F0FD", x"F406",
		x"F5FD", x"F6C8", x"F72A", x"F865", x"FB4A", x"0019", x"0637", x"0C5B",
		x"10D2", x"1232", x"101C", x"0B8B", x"069D", x"03A0", x"0417", x"0798",
		x"0CB4", x"112B", x"132D", x"11CC", x"0DD8", x"08D9", x"047C", x"01AB",
		x"008F", x"014C", x"037F", x"06C0", x"0AA4", x"0E8D", x"11CF", x"1357",
		x"1201", x"0DA1", x"06D2", x"FF03", x"F7C2", x"F24A", x"EF56", x"EF49",
		x"F1F9", x"F722", x"FE25", x"05EA", x"0CF6", x"11F0", x"1400", x"1314",
		x"1036", x"0C83", x"090E", x"0662", x"04A3", x"03AA", x"0354", x"03C3",
		x"0516", x"074B", x"0A1C", x"0D15", x"0FBD", x"11BF", x"12CC", x"12BE",
		x"1116", x"0D63", x"07A7", x"0074", x"F8ED", x"F261", x"EE00", x"EC4A",
		x"ED30", x"EFF8", x"F383", x"F6FC", x"F9F8", x"FBFC", x"FCDE", x"FC42",
		x"FA38", x"F6C3", x"F2A0", x"EEC8", x"ED14", x"EE96", x"F2F1", x"F8C4",
		x"FE2A", x"019B", x"027B", x"00EE", x"FD9C", x"F964", x"F589", x"F247",
		x"F00F", x"EF6D", x"F064", x"F2E4", x"F65E", x"FA5E", x"FE2B", x"00FB",
		x"0223", x"0100", x"FD85", x"F859", x"F295", x"EE2F", x"EC95", x"EE2B",
		x"F23B", x"F7A3", x"FD26", x"01FE", x"058D", x"07EB", x"097C", x"0B00",
		x"0C93", x"0E68", x"1042", x"11E9", x"1351", x"143A", x"14E1", x"1530",
		x"152D", x"14D8", x"141C", x"1309", x"114C", x"0F06", x"0C56", x"09B9",
		x"0769", x"05BF", x"054E", x"0601", x"07E4", x"0A92", x"0D7A", x"1029",
		x"1253", x"1381", x"13C9", x"12CB", x"1053", x"0C5F", x"06DA", x"FFCA",
		x"F82F", x"F15D", x"ED43", x"ECFD", x"F0E7", x"F82A", x"00F4", x"094B",
		x"0F78", x"1328", x"14F7", x"1590", x"1590", x"14C7", x"1284", x"0E0D",
		x"0731", x"FEBE", x"F687", x"F024", x"EC74", x"EB20", x"EB48", x"EBB4",
		x"EC1C", x"EC72", x"ED34", x"EE57", x"F007", x"F289", x"F5A4", x"F9BC",
		x"FE27", x"021D", x"04EB", x"05CA", x"046C", x"00C9", x"FB3C", x"F4E7",
		x"EF82", x"EC9F", x"ECEE", x"EFA5", x"F387", x"F753", x"F9E2", x"FAA8",
		x"F9B8", x"F767", x"F459", x"F10B", x"EDFB", x"EC06", x"EC3E", x"EF74",
		x"F582", x"FD6C", x"056A", x"0C41", x"1112", x"1393", x"135D", x"1081",
		x"0B05", x"038F", x"FB36", x"F3A0", x"EE2D", x"EB56", x"EA8C", x"EAB5",
		x"EADE", x"EACB", x"EB3A", x"EC68", x"EE1D", x"EFC1", x"F0CD", x"F114",
		x"F0B9", x"EFF0", x"EEED", x"EDB2", x"EC83", x"EBAD", x"EBCF", x"ED81",
		x"F118", x"F69F", x"FDAD", x"0557", x"0C48", x"1147", x"13CF", x"1435",
		x"1335", x"1158", x"0F0E", x"0CB7", x"0ABF", x"0963", x"08A3", x"08B3",
		x"0959", x"0ACF", x"0CED", x"0F6A", x"1193", x"131D", x"142B", x"14C4",
		x"151D", x"14C5", x"137A", x"10DA", x"0D6D", x"0A1F", x"0811", x"0825",
		x"0A3E", x"0DA1", x"10C1", x"1211", x"106A", x"0BAE", x"0557", x"FF9A",
		x"FC7F", x"FD1A", x"012E", x"0772", x"0DAA", x"11FA", x"12FD", x"10C5",
		x"0C5D", x"06E5", x"0193", x"FD07", x"F99F", x"F74C", x"F5FE", x"F547",
		x"F4E5", x"F4E6", x"F592", x"F6EF", x"F8C0", x"FAF9", x"FDB8", x"00FC",
		x"0482", x"07F1", x"0B13", x"0DCE", x"1001", x"11B7", x"1325", x"1420",
		x"14A8", x"14E4", x"149E", x"13EB", x"12BE", x"10F8", x"0E97", x"0C1D",
		x"0A55", x"0A1F", x"0BED", x"0F06", x"1210", x"1346", x"1193", x"0CB8",
		x"05EF", x"FF09", x"F9E0", x"F790", x"F83E", x"FB3A", x"FF80", x"0414",
		x"07F2", x"0A2F", x"0A55", x"07DC", x"0309", x"FC79", x"F579", x"EFC0",
		x"ECAE", x"ECC7", x"EF85", x"F3F1", x"F898", x"FC50", x"FEF9", x"00E5",
		x"0286", x"0451", x"064E", x"0895", x"0B06", x"0D86", x"0FFE", x"121E",
		x"13CF", x"14C4", x"1526", x"1534", x"1525", x"14EF", x"1458", x"1372",
		x"121A", x"105E", x"0E23", x"0BA3", x"0946", x"072F", x"0547", x"035B",
		x"015E", x"FEE8", x"FC01", x"F86C", x"F44F", x"F048", x"ED10", x"EB97",
		x"EC6A", x"EFC3", x"F587", x"FD2F", x"0584", x"0CE1", x"11F0", x"13C1",
		x"1233", x"0DDB", x"07EC", x"01CB", x"FCAB", x"F91A", x"F726", x"F6AA",
		x"F780", x"F999", x"FCD7", x"00F5", x"05E1", x"0AF5", x"0FB1", x"1300",
		x"143F", x"130D", x"0F9D", x"09FE", x"0292", x"FA56", x"F2D7", x"EDE8",
		x"ECDB", x"EFEC", x"F5C3", x"FCC4", x"02D9", x"069F", x"071B", x"03F6",
		x"FE29", x"F731", x"F125", x"EDC5", x"ED51", x"EF13", x"F17E", x"F315",
		x"F2FB", x"F15E", x"EEF2", x"ECAA", x"EB35", x"EA8E", x"EA55", x"EABC",
		x"EC4A", x"EF9B", x"F515", x"FC35", x"043F", x"0BB2", x"111D", x"134C",
		x"1195", x"0C8F", x"0547", x"FD68", x"F63C", x"F0BC", x"ED42", x"EB9A",
		x"EB30", x"EB22", x"EB53", x"EBD0", x"ECF5", x"EF1E", x"F1FE", x"F55E",
		x"F8F9", x"FCB5", x"0047", x"035A", x"05E3", x"07C0", x"0918", x"0A10",
		x"0A77", x"0A6D", x"0A02", x"0903", x"075A", x"04C7", x"011F", x"FC8A",
		x"F751", x"F239", x"EE51", x"ECA4", x"EE01", x"F262", x"F8EB", x"FFA5",
		x"04B4", x"072B", x"06DF", x"0458", x"0065", x"FBAE", x"F781", x"F480",
		x"F38D", x"F542", x"F98F", x"003B", x"07CD", x"0E99", x"129E", x"13A9",
		x"1292", x"1052", x"0E59", x"0D4D", x"0D86", x"0EB8", x"1098", x"1288",
		x"13FC", x"146F", x"12C2", x"0E88", x"07EB", x"0030", x"F89E", x"F24E",
		x"EDC3", x"EB2E", x"EA48", x"EA6E", x"EAD1", x"EB15", x"EB73", x"EC57",
		x"EDD7", x"EFE3", x"F260", x"F4F6", x"F78D", x"F9DD", x"FC39", x"FE99",
		x"0109", x"0389", x"05F6", x"0836", x"0A44", x"0C11", x"0DB9", x"0F3C",
		x"10C2", x"1244", x"13B8", x"1486", x"13E2", x"110E", x"0BAF", x"0460",
		x"FC31", x"F49B", x"EED1", x"EB59", x"EA1D", x"EA39", x"EADF", x"EB4B",
		x"EBAB", x"EC2B", x"ED77", x"F03C", x"F50C", x"FC14", x"047E", x"0C75",
		x"11F0", x"1456", x"141D", x"12F9", x"124C", x"12AF", x"13AD", x"140F",
		x"1257", x"0D6E", x"05BA", x"FC98", x"F41C", x"EE71", x"ECB9", x"EF10",
		x"F49C", x"FB82", x"01FE", x"06DD", x"099D", x"09C2", x"078C", x"0326",
		x"FD05", x"F640", x"F04D", x"ECFB", x"EDB4", x"F2BD", x"FA9E", x"033B",
		x"0AE9", x"1073", x"13C1", x"14BB", x"13C9", x"112C", x"0D7B", x"08FC",
		x"0438", x"FFD8", x"FC93", x"FADB", x"FB16", x"FCFC", x"008F", x"0599",
		x"0B43", x"102D", x"1303", x"12C7", x"0F93", x"0AA5", x"0526", x"0042",
		x"FCA4", x"FA33", x"F871", x"F6E9", x"F52D", x"F2E7", x"F061", x"EDF5",
		x"EC22", x"EC2F", x"EEA4", x"F3CD", x"FB25", x"0356", x"0AE7", x"1087",
		x"135D", x"129B", x"0EBE", x"08BC", x"01F0", x"FB98", x"F673", x"F2BC",
		x"F0A5", x"F01D", x"F121", x"F34D", x"F6AC", x"FAF6", x"0028", x"05A0",
		x"0AD7", x"0F47", x"1279", x"13D5", x"12E9", x"0F46", x"0927", x"0162",
		x"F954", x"F271", x"EDAB", x"EB7F", x"EBEA", x"EED7", x"F418", x"FB23",
		x"0307", x"0A74", x"1004", x"12CB", x"1212", x"0E29", x"0893", x"0377",
		x"0048", x"FFA0", x"00E1", x"039A", x"06F4", x"0A75", x"0D46", x"0EFC",
		x"0F20", x"0D71", x"09E1", x"047C", x"FDFC", x"F70B", x"F0FE", x"ED76",
		x"ED79", x"F1AB", x"F8F3", x"01BF", x"0A1E", x"1073", x"13EC", x"14D5",
		x"145D", x"13B4", x"13C0", x"1414", x"138C", x"10E0", x"0B4E", x"0392",
		x"FB34", x"F3EE", x"EED1", x"EBF9", x"EACA", x"EA7E", x"EAB5", x"EAEF",
		x"EB1F", x"EB3E", x"EB48", x"EB44", x"EB27", x"EB0A", x"EAF5", x"EAF1",
		x"EB30", x"EC60", x"EF2B", x"F42E", x"FB14", x"0310", x"0A7C", x"103F",
		x"1379", x"1486", x"140B", x"12EB", x"1208", x"11BF", x"1250", x"134F",
		x"1484", x"14FB", x"13FC", x"10FC", x"0B95", x"0448", x"FC22", x"F4A0",
		x"EF01", x"EC0E", x"EB5F", x"EBCC", x"EC42", x"EC16", x"EBA8", x"EB5E",
		x"EBBC", x"EC63", x"ECDF", x"ECCF", x"EC48", x"EBF7", x"ED3B", x"F0EE",
		x"F727", x"FECE", x"0664", x"0C79", x"1066", x"1210", x"123D", x"1161",
		x"0FA5", x"0D08", x"0933", x"043C", x"FE6A", x"F864", x"F2D5", x"EE78",
		x"EC4C", x"ECBF", x"EFF6", x"F534", x"FB3B", x"00E8", x"058C", x"091D",
		x"0B87", x"0D3C", x"0E7E", x"0F95", x"10C9", x"1223", x"1362", x"1447",
		x"14C9", x"14DD", x"149E", x"142E", x"1373", x"1287", x"1170", x"1034",
		x"0ED3", x"0D45", x"0B3E", x"0889", x"0539", x"0106", x"FC0B", x"F6C5",
		x"F19A", x"EDA6", x"EC0C", x"ED6A", x"F1FB", x"F8C2", x"0096", x"0811",
		x"0E18", x"1256", x"1434", x"13B7", x"1097", x"0AF1", x"034B", x"FAE0",
		x"F371", x"EE83", x"ED13", x"EEC0", x"F272", x"F67B", x"F910", x"F924",
		x"F6C3", x"F2E4", x"EF01", x"ECB7", x"ED66", x"F19A", x"F8F6", x"0228",
		x"0AD9", x"110E", x"133B", x"1168", x"0CD5", x"07C0", x"0407", x"02EB",
		x"04E0", x"093E", x"0E6C", x"1225", x"12A3", x"0FC9", x"0B7D", x"07BA",
		x"06A0", x"08AB", x"0CB6", x"10BD", x"125B", x"1051", x"0B0D", x"0434",
		x"FDC6", x"F8BD", x"F5A7", x"F3E5", x"F312", x"F272", x"F152", x"EF79",
		x"ED61", x"EC42", x"ED10", x"F050", x"F631", x"FD91", x"0558", x"0BEA",
		x"109F", x"1336", x"1475", x"14B5", x"1468", x"13D6", x"133D", x"128C",
		x"11BC", x"107F", x"0EFC", x"0D6C", x"0C02", x"0AA5", x"08E7", x"061F",
		x"01FE", x"FC91", x"F6A1", x"F12E", x"EDA5", x"ED20", x"EFB1", x"F480",
		x"F9FC", x"FDEF", x"FED7", x"FC82", x"F7BD", x"F26E", x"EE87", x"ED79",
		x"F050", x"F67E", x"FE9F", x"06EA", x"0DA7", x"1217", x"142A", x"1424",
		x"11DC", x"0D2F", x"062C", x"FDA3", x"F553", x"EF3E", x"ECB6", x"EDD2",
		x"F141", x"F4E2", x"F6D4", x"F614", x"F306", x"EF4A", x"ECE4", x"ED68",
		x"F15C", x"F767", x"FDBD", x"022D", x"03B1", x"0248", x"FF02", x"FB00",
		x"F70A", x"F3CB", x"F1EB", x"F1D6", x"F414", x"F8B1", x"FF15", x"0687",
		x"0D43", x"11CF", x"130E", x"10AD", x"0B51", x"03E8", x"FBFE", x"F4CE",
		x"EF97", x"EC95", x"EBF2", x"ED63", x"F03B", x"F38E", x"F6B5", x"F976",
		x"FBAE", x"FDB4", x"FF92", x"0189", x"03DE", x"06AA", x"09AB", x"0C9F",
		x"0F3B", x"1160", x"12D2", x"13A8", x"13F1", x"13D3", x"138C", x"1328",
		x"1287", x"118D", x"0FE6", x"0D08", x"08B5", x"02CF", x"FBE4", x"F4D1",
		x"EF2B", x"ECA7", x"EDA3", x"F0DA", x"F456", x"F5D1", x"F4B2", x"F1B8",
		x"EED7", x"EE1A", x"F0A8", x"F64D", x"FCC7", x"0180", x"023B", x"FED3",
		x"F8CE", x"F277", x"EE35", x"ED33", x"EF39", x"F32C", x"F72A", x"F9BA",
		x"FA45", x"F915", x"F6A5", x"F38F", x"F055", x"ED66", x"EBB4", x"EBE5",
		x"EEAD", x"F406", x"FB6A", x"036F", x"0AD9", x"103A", x"135D", x"1493",
		x"14A2", x"13E6", x"1290", x"1088", x"0DF0", x"0B37", x"0917", x"0800",
		x"0808", x"0907", x"0AD7", x"0D15", x"0F51", x"114A", x"12E1", x"13F4",
		x"1486", x"148E", x"13D8", x"1275", x"10C8", x"0F4A", x"0E70", x"0EED",
		x"109E", x"12A9", x"13D7", x"12EA", x"0F26", x"08DE", x"0110", x"F975",
		x"F335", x"EF01", x"EC81", x"EB5E", x"EB0B", x"EB12", x"EB07", x"EAFB",
		x"EB07", x"EB95", x"ED1F", x"EF76", x"F206", x"F491", x"F686", x"F72A",
		x"F614", x"F369", x"EFE8", x"ECF6", x"EBE4", x"ED68", x"F1AB", x"F7FE",
		x"FF49", x"0666", x"0C4B", x"1090", x"130D", x"1449", x"14C8", x"14C8",
		x"1491", x"13F2", x"127B", x"0FA1", x"0B18", x"04A7", x"FD0B", x"F5C1",
		x"EFFB", x"ECDB", x"ED69", x"F1AF", x"F8F2", x"017A", x"0938", x"0F1B",
		x"12A8", x"145E", x"14F8", x"1504", x"14BC", x"1437", x"1319", x"1167",
		x"0F7C", x"0E3E", x"0E53", x"0FEA", x"1234", x"13AB", x"129A", x"0E2F",
		x"0735", x"FF04", x"F7B2", x"F271", x"EF6C", x"EDFE", x"ED64", x"ECFA",
		x"EC5E", x"EBB4", x"EB3C", x"EBB7", x"EE51", x"F38B", x"FAE6", x"0312",
		x"0A72", x"1018", x"13A2", x"1561", x"15BF", x"1560", x"14CC", x"13E4",
		x"1287", x"10B2", x"0EC8", x"0D22", x"0C1C", x"0BDD", x"0C92", x"0E2C",
		x"1039", x"124B", x"13CE", x"14B2", x"146B", x"12CC", x"0F46", x"09DD",
		x"02BE", x"FACE", x"F381", x"EE36", x"EC1D", x"ED64", x"F174", x"F7D1",
		x"FF4F", x"06D3", x"0D20", x"1194", x"1403", x"14CE", x"148E", x"13A0",
		x"127E", x"10FC", x"0F94", x"0E35", x"0CA7", x"0AB3", x"07E8", x"0444",
		x"0022", x"FC01", x"F888", x"F624", x"F594", x"F753", x"FBCF", x"0283",
		x"09F0", x"0FCD", x"129F", x"1250", x"103E", x"0E53", x"0E19", x"0FA4",
		x"11C2", x"1237", x"0F14", x"089B", x"00B2", x"FA98", x"F89F", x"FB8F",
		x"023D", x"09F1", x"0FF4", x"1273", x"11AB", x"0F78", x"0D9D", x"0DA3",
		x"0F74", x"11CA", x"1262", x"0F8C", x"0939", x"0175", x"FAE6", x"F731",
		x"F67A", x"F81A", x"FB6B", x"FFC1", x"042C", x"07E1", x"0A38", x"0AE7",
		x"0A21", x"0824", x"054D", x"020C", x"FEBA", x"FBBD", x"F979", x"F852",
		x"F84D", x"F952", x"FB68", x"FE23", x"0163", x"04B5", x"0800", x"0AF7",
		x"0D8D", x"0FA3", x"115C", x"129E", x"1391", x"146D", x"14E6", x"151B",
		x"150D", x"1480", x"1359", x"1196", x"0F70", x"0D08", x"0B35", x"0A46",
		x"0A36", x"0AE6", x"0C45", x"0E02", x"0FC8", x"1171", x"12C2", x"13B5",
		x"1457", x"14A2", x"149C", x"144B", x"13C6", x"12BC", x"10D9", x"0DEC",
		x"09F7", x"0514", x"FF2C", x"F8BD", x"F2C5", x"EE4C", x"EC2B", x"ECE3",
		x"F0B4", x"F70C", x"FF03", x"0717", x"0DD4", x"1245", x"13E5", x"12E1",
		x"0FEC", x"0BB2", x"0711", x"02C7", x"FF17", x"FC06", x"F983", x"F745",
		x"F526", x"F350", x"F1B1", x"F049", x"EF2E", x"EE6C", x"EDC5", x"ED2E",
		x"EC30", x"EB74", x"EBDE", x"EE62", x"F3B5", x"FB83", x"0438", x"0BFF",
		x"11A1", x"14ED", x"164D", x"1603", x"13DC", x"0F79", x"0918", x"0142",
		x"F90F", x"F198", x"EC8C", x"EAF2", x"ED50", x"F2DF", x"FAB6", x"032D",
		x"0AC7", x"10BA", x"148D", x"1627", x"1561", x"1261", x"0D37", x"064F",
		x"FE52", x"F65C", x"EFC0", x"EC09", x"EB9E", x"EE8A", x"F450", x"FBDE",
		x"043D", x"0BD4", x"1190", x"149B", x"157C", x"1540", x"14D3", x"1479",
		x"13FA", x"1327", x"11DC", x"1098", x"0FBC", x"0F96", x"1049", x"11BC",
		x"1353", x"147C", x"1513", x"1518", x"149F", x"13C3", x"12C7", x"11A6",
		x"104B", x"0E78", x"0C65", x"0A17", x"07BF", x"0522", x"025A", x"FFAC",
		x"FD40", x"FAF5", x"F88D", x"F5EC", x"F361", x"F129", x"EF5D", x"EDCA",
		x"EC6B", x"EB75", x"EAEF", x"EAF5", x"EB20", x"EB1F", x"EAF1", x"EAD7",
		x"EB09", x"EBA4", x"EC94", x"EDC3", x"EEED", x"EF65", x"EEE3", x"ED6B",
		x"EC2F", x"EC84", x"EF7C", x"F585", x"FD79", x"05F3", x"0D14", x"11D9",
		x"13C9", x"12E9", x"0F77", x"0A02", x"032C", x"FBA4", x"F49F", x"EF52",
		x"EC92", x"ECE8", x"F042", x"F5FC", x"FCF1", x"03FE", x"0A3E", x"0EF9",
		x"1225", x"13F4", x"14C6", x"1504", x"1506", x"14D7", x"1487", x"13D9",
		x"12AB", x"10D5", x"0E2A", x"0AD8", x"0758", x"04B4", x"03DA", x"054F",
		x"08C7", x"0D1F", x"10EA", x"12B5", x"1181", x"0D66", x"07E4", x"033A",
		x"0126", x"0266", x"0659", x"0B49", x"0FC0", x"1222", x"1149", x"0CB6",
		x"04FD", x"FBD0", x"F39D", x"EE51", x"ECA9", x"EE25", x"F19C", x"F536",
		x"F778", x"F74B", x"F481", x"F06F", x"ED52", x"ED3E", x"F09C", x"F675",
		x"FCA6", x"013C", x"0336", x"0268", x"FF8A", x"FB5E", x"F6D8", x"F2EE",
		x"F014", x"EEC7", x"EF37", x"F12D", x"F47A", x"F855", x"FC64", x"FF95",
		x"012C", x"009C", x"FDBB", x"F936", x"F3C0", x"EF08", x"EC7C", x"ED0A",
		x"F090", x"F616", x"FC35", x"01B2", x"0613", x"092C", x"0B46", x"0CBC",
		x"0DFD", x"0F4E", x"10B9", x"1239", x"1389", x"145B", x"14C3", x"14BB",
		x"145E", x"141D", x"13E2", x"13D5", x"13FC", x"143E", x"1456", x"140A",
		x"135B", x"12AC", x"1220", x"1231", x"12DA", x"13CE", x"1482", x"14D0",
		x"14BA", x"1451", x"142D", x"143A", x"145F", x"1413", x"1282", x"0EDF",
		x"089B", x"0062", x"F7B4", x"F08C", x"EC7B", x"EC28", x"EF7D", x"F5A7",
		x"FD13", x"044D", x"09FD", x"0DE0", x"1040", x"1170", x"11D9", x"1109",
		x"0F28", x"0C37", x"0895", x"048B", x"0075", x"FCD3", x"F9F2", x"F788",
		x"F5AF", x"F3FB", x"F288", x"F12B", x"EFAB", x"EE10", x"EC77", x"EB89",
		x"EB61", x"EBF3", x"ECC3", x"ED17", x"ECC4", x"EBED", x"EB7C", x"EC83",
		x"F004", x"F60E", x"FDED", x"0607", x"0CC7", x"10E0", x"124D", x"1166",
		x"0EDD", x"0B22", x"06D4", x"02E9", x"0063", x"006B", x"0313", x"0809",
		x"0DAA", x"11B4", x"1284", x"0FAE", x"0B03", x"06DD", x"0523", x"0692",
		x"0A85", x"0F10", x"1211", x"11CC", x"0E50", x"086C", x"01C5", x"FB68",
		x"F648", x"F2B7", x"F086", x"EF4F", x"EE7E", x"EE0C", x"EDD1", x"EDF0",
		x"EE52", x"EF55", x"F0F7", x"F332", x"F5D6", x"F8C1", x"FBD5", x"FF1A",
		x"0250", x"0529", x"079E", x"09A1", x"0B44", x"0CDF", x"0E86", x"1039",
		x"11F4", x"136C", x"1471", x"14B5", x"1441", x"138B", x"1329", x"13A8",
		x"142C", x"139B", x"1108", x"0BE7", x"04D2", x"FCC2", x"F56E", x"F02E",
		x"ED71", x"ECF6", x"EE13", x"F044", x"F334", x"F65F", x"F958", x"FB0B",
		x"FACE", x"F869", x"F46B", x"F025", x"ED25", x"ECD9", x"EFE0", x"F5E4",
		x"FDE1", x"0620", x"0D53", x"1229", x"141F", x"1302", x"0F65", x"09FC",
		x"03E4", x"FDFC", x"F8BA", x"F477", x"F16D", x"EF5C", x"EE16", x"ED67",
		x"ED2C", x"ED28", x"ED60", x"EDE0", x"EEEB", x"F079", x"F2CE", x"F590",
		x"F8B3", x"FBB6", x"FE73", x"00AE", x"0292", x"0435", x"05DC", x"07C5",
		x"0A73", x"0DA9", x"1100", x"1326", x"12DE", x"0F79", x"0949", x"01D6",
		x"FA9D", x"F549", x"F2E5", x"F436", x"F90A", x"004D", x"0801", x"0E45",
		x"1206", x"133D", x"128C", x"116B", x"111D", x"11E6", x"132F", x"1439",
		x"1495", x"1489", x"1492", x"14CB", x"148D", x"133C", x"0FEC", x"0A84",
		x"0320", x"FAD6", x"F315", x"EDCD", x"EC37", x"EE8C", x"F3E4", x"FAFD",
		x"027D", x"095C", x"0ECD", x"122F", x"13C0", x"13D2", x"12CF", x"10F0",
		x"0E7A", x"0B8D", x"08C4", x"06BB", x"05E1", x"0645", x"07DE", x"0A4D",
		x"0CFE", x"0F7E", x"1179", x"12BE", x"135D", x"1384", x"1346", x"12DF",
		x"121A", x"10BE", x"0E96", x"0B3D", x"0695", x"009C", x"F9CA", x"F339",
		x"EE5D", x"EC5B", x"ED67", x"F0A7", x"F4BC", x"F7DA", x"F924", x"F83B",
		x"F5DA", x"F2C9", x"EFF3", x"EDCC", x"EC70", x"EBCB", x"EBDC", x"EC9E",
		x"EDDB", x"EFC4", x"F20E", x"F47F", x"F668", x"F7B4", x"F844", x"F845",
		x"F7B5", x"F682", x"F48F", x"F1F7", x"EF3A", x"ECBF", x"EB81", x"EC32",
		x"EF9F", x"F56D", x"FCDA", x"047B", x"0B2B", x"1046", x"134F", x"1495",
		x"14AA", x"1404", x"12DC", x"1115", x"0E9D", x"0B89", x"0811", x"0453",
		x"00A4", x"FD77", x"FACC", x"F8A8", x"F6C1", x"F552", x"F42E", x"F3A9",
		x"F38D", x"F3E9", x"F4B4", x"F63B", x"F8A9", x"FC51", x"0141", x"06F7",
		x"0CAE", x"1130", x"135C", x"12B0", x"0F3F", x"0A06", x"0425", x"FECA",
		x"FADF", x"F898", x"F810", x"F8FD", x"FB58", x"FF18", x"03FE", x"0985",
		x"0EA9", x"1263", x"1391", x"11DB", x"0D75", x"077C", x"012E", x"FBA2",
		x"F744", x"F44F", x"F300", x"F2FC", x"F42F", x"F690", x"FAAB", x"00DD",
		x"0807", x"0D7A", x"0E91", x"0B3F", x"0657", x"0422", x"0693", x"0C3C",
		x"11D3", x"151E", x"1601", x"1590", x"14F7", x"140E", x"12AF", x"103C",
		x"0C8B", x"078A", x"012D", x"FA32", x"F3BE", x"EEE7", x"EC64", x"EC74",
		x"EF06", x"F33D", x"F806", x"FC47", x"FF80", x"01A8", x"0349", x"04E2",
		x"06DA", x"099C", x"0D3F", x"10EC", x"1388", x"1391", x"102B", x"0A0C",
		x"0292", x"FB58", x"F59A", x"F1AB", x"EF68", x"EE25", x"ED38", x"EC5B",
		x"EB8E", x"EAD9", x"EADD", x"EC12", x"EEEA", x"F395", x"F9F7", x"016A",
		x"08DD", x"0F31", x"133A", x"1434", x"1210", x"0D0E", x"064E", x"FEEE",
		x"F7E3", x"F204", x"EDBF", x"EBC0", x"ECB3", x"F096", x"F6B4", x"FDFE",
		x"057C", x"0C56", x"118A", x"1446", x"1409", x"10FC", x"0BA3", x"04CC",
		x"FD3F", x"F615", x"F066", x"ED08", x"EC69", x"EE5B", x"F297", x"F88D",
		x"FF6C", x"066D", x"0CB1", x"1145", x"134B", x"1203", x"0D11", x"0577",
		x"FCC2", x"F52E", x"EFA7", x"EC77", x"EB0F", x"EB01", x"EC7C", x"EFD5",
		x"F54F", x"FC96", x"04E8", x"0C74", x"11D0", x"1385", x"116B", x"0C6A",
		x"05D3", x"FEAB", x"F7C4", x"F1DE", x"EDC0", x"EC06", x"ECD9", x"F037",
		x"F5E7", x"FD30", x"04E6", x"0BDA", x"10E1", x"1380", x"1368", x"1094",
		x"0B88", x"04E8", x"FD89", x"F6AB", x"F0F7", x"ED21", x"EC3D", x"EF12",
		x"F5A0", x"FE61", x"0715", x"0E12", x"12B0", x"1539", x"15BD", x"147F",
		x"1128", x"0BB6", x"046F", x"FC6F", x"F4D7", x"EF19", x"EBCB", x"EADD",
		x"EC23", x"EF9C", x"F551", x"FCEF", x"05AB", x"0D8B", x"1295", x"13A5",
		x"110C", x"0C12", x"059D", x"FE9D", x"F7A2", x"F1A5", x"ED9A", x"EC3D",
		x"EDEE", x"F27C", x"F931", x"00F2", x"0850", x"0E44", x"127B", x"14A1",
		x"1503", x"1440", x"12A3", x"10DA", x"0EFD", x"0D2B", x"0B99", x"0A29",
		x"08AD", x"06DA", x"04F0", x"02E3", x"00B3", x"FE04", x"FAAB", x"F6DA",
		x"F2FA", x"EF83", x"ED04", x"EC0F", x"ED67", x"F17E", x"F801", x"0003",
		x"080F", x"0EB7", x"12DF", x"1446", x"12DB", x"0F1C", x"0992", x"0292",
		x"FB0B", x"F402", x"EF2D", x"ED95", x"EFDF", x"F547", x"FC1D", x"02E6",
		x"07B8", x"0954", x"0719", x"0152", x"F9A4", x"F282", x"EE18", x"ECE0",
		x"EDD4", x"EF25", x"EF71", x"EEA5", x"EDD0", x"EEDA", x"F31D", x"FA44",
		x"0286", x"08CF", x"0AE7", x"081B", x"016E", x"F933", x"F204", x"EDD4",
		x"ECBB", x"EDA4", x"EEB8", x"EEBB", x"EDA6", x"ECCF", x"EDDB", x"F1FB",
		x"F8E0", x"00F6", x"086D", x"0DEE", x"1170", x"137F", x"149D", x"151E",
		x"154D", x"1551", x"1530", x"1506", x"1484", x"136E", x"11FD", x"1030",
		x"0E16", x"0BD4", x"0992", x"073C", x"04D9", x"0279", x"FFE9", x"FD10",
		x"FA15", x"F738", x"F49D", x"F258", x"F074", x"EEF4", x"EDCC", x"ECFA",
		x"EC54", x"EBCE", x"EB41", x"EB45", x"ECAA", x"F091", x"F737", x"FFA8",
		x"0806", x"0EA4", x"12DB", x"150F", x"15C2", x"150D", x"1275", x"0E1F",
		x"07CA", x"000B", x"F814", x"F16D", x"ED3C", x"EC0A", x"ED88", x"F190",
		x"F7E5", x"0005", x"088D", x"0F7D", x"1335", x"1304", x"0F3D", x"0920",
		x"020C", x"FB0A", x"F4C8", x"EFD2", x"ECE5", x"EC95", x"EFA5", x"F5E3",
		x"FE24", x"06AC", x"0DA8", x"123A", x"1496", x"154D", x"153A", x"14E6",
		x"14E6", x"14E4", x"1496", x"13CD", x"12CD", x"11B1", x"10C4", x"103D",
		x"1043", x"1138", x"1268", x"13AA", x"144F", x"141D", x"12AF", x"0FD6",
		x"0B78", x"05B2", x"FEC6", x"F7B7", x"F176", x"ED72", x"EC74", x"EECB",
		x"F40F", x"FB51", x"0358", x"0A83", x"1001", x"133E", x"147F", x"140D",
		x"1243", x"0FB8", x"0CAC", x"09C8", x"0747", x"0599", x"04E3", x"0527",
		x"0674", x"08CD", x"0BBB", x"0ED2", x"1168", x"133D", x"143D", x"13F7",
		x"11B9", x"0CF2", x"05A7", x"FD73", x"F5C0", x"EFD3", x"EC0D", x"EA2F",
		x"E9D6", x"EABA", x"ED79", x"F23F", x"F925", x"0152", x"095D", x"0FC8",
		x"12F2", x"1261", x"0E1A", x"070B", x"FEB6", x"F6AD", x"F03A", x"EC1B",
		x"EA8D", x"EA9E", x"EB53", x"EB9B", x"EB8F", x"EB8D", x"EBF2", x"ECDA",
		x"EDD9", x"EE6E", x"EE45", x"ED73", x"EC81", x"EBB9", x"EB5C", x"EB4F",
		x"EB74", x"EB8F", x"EB5B", x"EB0C", x"EABC", x"EABA", x"EB49", x"EC47",
		x"ED73", x"EE2E", x"EE71", x"EDE2", x"ED0A", x"EC2E", x"EB87", x"EB52",
		x"EB70", x"EC07", x"ED31", x"EEDD", x"F0FB", x"F355", x"F5CF", x"F826",
		x"FA2E", x"FB87", x"FBFF", x"FB76", x"FA09", x"F7B1", x"F4D9", x"F234",
		x"EFF6", x"EE6F", x"ED8D", x"ED08", x"ED41", x"EE41", x"F015", x"F295",
		x"F585", x"F8C9", x"FC19", x"FF1C", x"01A5", x"03CD", x"0572", x"06CD",
		x"086D", x"0AB8", x"0DD6", x"1119", x"133E", x"1379", x"116A", x"0D0C",
		x"06D8", x"FF82", x"F853", x"F24C", x"EE09", x"EBB4", x"EAAA", x"EA8C",
		x"EAE9", x"EB78", x"EC34", x"ECE1", x"ED6A", x"EE0E", x"EEEB", x"F02F",
		x"F1E8", x"F459", x"F789", x"FB69", x"FFFE", x"050C", x"0A51", x"0F40",
		x"12E5", x"1406", x"1204", x"0CF5", x"056B", x"FCCA", x"F4AD", x"EEEE",
		x"ECAC", x"EDFC", x"F1B3", x"F5DD", x"F8C3", x"F996", x"F808", x"F4B3",
		x"F0A1", x"ED53", x"EC59", x"EF09", x"F529", x"FDAA", x"06C0", x"0E67",
		x"12CC", x"134A", x"1057", x"0B7D", x"0718", x"04BB", x"059C", x"092F",
		x"0DF3", x"118A", x"1215", x"0F47", x"0A4C", x"05A9", x"03B8", x"054D",
		x"09BF", x"0EC3", x"11F3", x"11EC", x"0EB6", x"0996", x"0467", x"00A2",
		x"FF20", x"FFD5", x"0256", x"05C9", x"09B3", x"0D9C", x"1101", x"133A",
		x"1378", x"1189", x"0D2F", x"06DF", x"FF70", x"F83E", x"F243", x"EE1F",
		x"EBCF", x"EABB", x"EA93", x"EAE0", x"EB59", x"EBF6", x"ECB6", x"EDB2",
		x"EF05", x"F090", x"F278", x"F492", x"F6D1", x"F933", x"FBC4", x"FEF1",
		x"026B", x"0655", x"0A06", x"0D47", x"0FB3", x"114E", x"122C", x"1203",
		x"10BC", x"0E0A", x"099D", x"036A", x"FC06", x"F4A7", x"EF01", x"EC60",
		x"ED73", x"F1BD", x"F80E", x"FF1E", x"0624", x"0C47", x"10FB", x"138D",
		x"1369", x"0FF6", x"0981", x"00E9", x"F7FF", x"F0C3", x"EC76", x"EACC",
		x"EAC8", x"EB20", x"EB74", x"EC72", x"EF28", x"F45B", x"FBA5", x"03E4",
		x"0B6C", x"10EA", x"1402", x"14D4", x"1415", x"127B", x"10EC", x"1005",
		x"103F", x"116A", x"12EB", x"138B", x"1234", x"0E48", x"07ED", x"004D",
		x"F911", x"F3DC", x"F1C1", x"F33C", x"F7E4", x"FEDE", x"0688", x"0D58",
		x"11D8", x"132A", x"1183", x"0E46", x"0B15", x"08EA", x"0802", x"0786",
		x"063A", x"037D", x"FF06", x"F96B", x"F3BC", x"EF55", x"ED34", x"EE0A",
		x"F19D", x"F6F6", x"FC44", x"001F", x"01CB", x"018F", x"FFFE", x"FD81",
		x"FA5B", x"F6A4", x"F2EF", x"EFC7", x"ED5D", x"EBDA", x"EB2F", x"EB38",
		x"EBB9", x"EC21", x"EC1B", x"EBB8", x"EBB2", x"ECFD", x"F08A", x"F643",
		x"FDAC", x"05A3", x"0C8A", x"1112", x"12A8", x"113E", x"0D17", x"06C0",
		x"FEE2", x"F6BC", x"F026", x"EC68", x"EBB7", x"ED38", x"EF6D", x"F131",
		x"F227", x"F2C7", x"F3F6", x"F660", x"FA60", x"FFFC", x"06AD", x"0D3B",
		x"11F0", x"138B", x"11DF", x"0E31", x"0A26", x"0730", x"0637", x"074E",
		x"09BF", x"0CD5", x"0FA7", x"11F6", x"1374", x"1432", x"13E0", x"129C",
		x"1077", x"0DA2", x"0A5F", x"072E", x"055A", x"05C7", x"08B4", x"0D1B",
		x"1115", x"12D1", x"113C", x"0C9D", x"0686", x"015C", x"FF2E", x"00D0",
		x"059A", x"0B99", x"1095", x"12CF", x"1189", x"0D68", x"07C6", x"0223",
		x"FD9E", x"FA71", x"F85D", x"F6FB", x"F5B7", x"F447", x"F28C", x"F0A5",
		x"EEB8", x"ECEB", x"EB9B", x"EAD0", x"EA90", x"EAB6", x"EB00", x"EB13",
		x"EB29", x"EB37", x"EB98", x"EC46", x"ED7D", x"EEC4", x"EFD4", x"F065",
		x"EFF3", x"EE9F", x"ED0F", x"EBD8", x"EB44", x"EB1D", x"EAF2", x"EAB3",
		x"EB0E", x"ED01", x"F157", x"F816", x"0038", x"085A", x"0EF5", x"12E2",
		x"13DD", x"11E5", x"0D42", x"0682", x"FE7C", x"F672", x"EFE1", x"EBAA",
		x"EA1C", x"EA50", x"EB19", x"EB82", x"EB82", x"EBC8", x"ECD8", x"EED3",
		x"F149", x"F3DA", x"F635", x"F869", x"FA9F", x"FCD5", x"FF26", x"019B",
		x"0451", x"0722", x"0A25", x"0CDB", x"0F4E", x"116A", x"1329", x"143D",
		x"14E1", x"1503", x"1487", x"13B5", x"124D", x"106F", x"0E1D", x"0BAC",
		x"0994", x"0836", x"0856", x"09E8", x"0CBC", x"0FC2", x"1247", x"13E5",
		x"14DB", x"151F", x"140B", x"1103", x"0BBD", x"0477", x"FC55", x"F4CE",
		x"EF29", x"EBD3", x"EAA8", x"EB2E", x"ED16", x"F0B3", x"F660", x"FE0E",
		x"0677", x"0DEA", x"12B5", x"1499", x"147B", x"1391", x"128A", x"11AC",
		x"10D7", x"0FEA", x"0EC8", x"0D08", x"0AA4", x"07F2", x"0510", x"0218",
		x"FF24", x"FC6D", x"F9FC", x"F7E9", x"F5DF", x"F399", x"F13C", x"EEEE",
		x"ECF8", x"EBA7", x"EADB", x"EA95", x"EABA", x"EB75", x"ECCF", x"EEFF",
		x"F1A9", x"F44F", x"F618", x"F616", x"F44B", x"F15B", x"EEC3", x"EE49",
		x"F0E1", x"F64F", x"FD2C", x"02F6", x"05A0", x"0422", x"FED8", x"F7A8",
		x"F118", x"ED72", x"ED0A", x"EEF6", x"F127", x"F1E6", x"F0C3", x"EE61",
		x"ECD6", x"EE33", x"F330", x"FACD", x"02DA", x"097A", x"0E20", x"10FB",
		x"128E", x"1364", x"13CF", x"1428", x"149F", x"14FE", x"1529", x"148C",
		x"1349", x"1192", x"0FD6", x"0E45", x"0D18", x"0C71", x"0C8F", x"0DB2",
		x"0F5B", x"1153", x"12F6", x"1410", x"14A0", x"14F8", x"1511", x"1529",
		x"153A", x"1511", x"14CE", x"1410", x"1269", x"0F66", x"0A71", x"0383",
		x"FB80", x"F40A", x"EECC", x"EC86", x"ED0E", x"EEDB", x"F054", x"F06C",
		x"EEE0", x"ECF4", x"EC93", x"EF40", x"F501", x"FC89", x"038F", x"0896",
		x"0AFA", x"0AFF", x"08F3", x"0530", x"008B", x"FBA1", x"F791", x"F486",
		x"F280", x"F104", x"EFF0", x"EF16", x"EE30", x"ED4C", x"EC3E", x"EBB4",
		x"EC8C", x"EFDF", x"F5DE", x"FD9D", x"0589", x"0C4C", x"1128", x"13F1",
		x"1519", x"154F", x"1509", x"1483", x"1365", x"11B7", x"0F92", x"0D9C",
		x"0C69", x"0C8B", x"0DD2", x"100C", x"1233", x"13D3", x"14BD", x"1544",
		x"159C", x"1509", x"1241", x"0CB5", x"04F6", x"FC6F", x"F4BE", x"EEFA",
		x"EBA3", x"EAC2", x"EC78", x"F089", x"F6C7", x"FE95", x"06C9", x"0DF9",
		x"1302", x"157F", x"161D", x"15DD", x"1573", x"1504", x"1423", x"1296",
		x"1058", x"0D7B", x"0A36", x"06D2", x"038E", x"0082", x"FDCA", x"FBBD",
		x"F9EB", x"F8CA", x"F87D", x"F942", x"FB33", x"FE39", x"01B9", x"0534",
		x"082A", x"0A57", x"0B5D", x"0AF7", x"0968", x"06D2", x"0383", x"FFE6",
		x"FCB3", x"FA1C", x"F8A0", x"F8CD", x"FAB6", x"FE14", x"023D", x"0664",
		x"09C9", x"0BDE", x"0C1A", x"09F3", x"054E", x"FEB1", x"F756", x"F0E7",
		x"ED07", x"EC3F", x"EDBA", x"F01E", x"F1F4", x"F286", x"F1B1", x"F01B",
		x"EE05", x"EC68", x"EB78", x"EB6A", x"EBF6", x"ECCD", x"EDD2", x"EF1F",
		x"F0A5", x"F273", x"F455", x"F66D", x"F8E7", x"FB82", x"FE18", x"0067",
		x"02A4", x"04EB", x"0786", x"0A29", x"0CA7", x"0F11", x"1143", x"130F",
		x"144C", x"1516", x"1576", x"15A2", x"15A0", x"1573", x"1557", x"1565",
		x"1550", x"1506", x"1450", x"12C7", x"0FEA", x"0B32", x"0479", x"FC93",
		x"F4EC", x"EF0B", x"EC0D", x"EBD4", x"ED13", x"EE4F", x"EE56", x"ED54",
		x"EC80", x"ED81", x"F187", x"F871", x"0131", x"09A5", x"1019", x"139A",
		x"13AD", x"10C3", x"0B8B", x"04F6", x"FE0A", x"F7E1", x"F334", x"EFF9",
		x"EDF6", x"ECA0", x"EBD4", x"EB31", x"EAD1", x"EAC5", x"EBB4", x"EE82",
		x"F3CF", x"FB2A", x"0374", x"0B09", x"10AB", x"13FE", x"1552", x"1593",
		x"156E", x"1535", x"1491", x"1388", x"121C", x"10ED", x"107A", x"10FF",
		x"125A", x"13AB", x"13C6", x"118D", x"0C88", x"050D", x"FC68", x"F46D",
		x"EEF1", x"ED4B", x"EFCD", x"F585", x"FCB8", x"0379", x"088E", x"0AFC",
		x"0A57", x"06C0", x"00D2", x"F9D5", x"F343", x"EE83", x"EC78", x"ED51",
		x"F064", x"F4A3", x"F8BC", x"FBFD", x"FE27", x"FF9C", x"00EB", x"0282",
		x"0474", x"0689", x"0895", x"0A63", x"0BED", x"0D80", x"0F57", x"1188",
		x"1391", x"1466", x"132F", x"0F48", x"0912", x"0189", x"F9EE", x"F3AA",
		x"EF4A", x"ECEB", x"EBEF", x"EBF3", x"EC49", x"ED22", x"EED6", x"F191",
		x"F5C0", x"FBA8", x"02CC", x"0A31", x"1045", x"1353", x"12AE", x"0F67",
		x"0B6D", x"08F6", x"0949", x"0C1F", x"0FEC", x"1268", x"11B2", x"0D77",
		x"074C", x"021A", x"FFF4", x"01DD", x"06ED", x"0CF2", x"117B", x"12E5",
		x"110A", x"0D07", x"0886", x"04F2", x"0319", x"0365", x"0587", x"08C5",
		x"0C8D", x"1022", x"12EF", x"148C", x"1406", x"1123", x"0BFF", x"052B",
		x"FDC6", x"F6D2", x"F129", x"ED87", x"EBC7", x"EB78", x"EC00", x"ECBC",
		x"ED8D", x"EE09", x"EE37", x"EE1D", x"EDE0", x"ED78", x"ECDE", x"EC16",
		x"EB4F", x"EAF2", x"EB23", x"EBFD", x"ED83", x"EFCE", x"F2B2", x"F5C7",
		x"F894", x"FA86", x"FB60", x"FB02", x"F923", x"F5E7", x"F207", x"EE9D",
		x"ECBD", x"EDAC", x"F177", x"F826", x"007F", x"08F1", x"0FA0", x"1361",
		x"1419", x"122E", x"0E7D", x"0974", x"03BF", x"FDCD", x"F85C", x"F3D4",
		x"F08C", x"EE2A", x"ECC5", x"EC5F", x"ECF8", x"EEE6", x"F292", x"F7FA",
		x"FEC7", x"0617", x"0CAB", x"1162", x"13A4", x"1396", x"116C", x"0DCE",
		x"0970", x"0532", x"01FB", x"0078", x"00F7", x"0374", x"078F", x"0C72",
		x"10C5", x"12FE", x"1229", x"0E57", x"090F", x"04B7", x"0350", x"0595",
		x"0A3F", x"0F69", x"12BA", x"12D8", x"0FD3", x"0AD2", x"0587", x"0198",
		x"FFE5", x"0072", x"02F0", x"06C5", x"0B1B", x"0F37", x"127E", x"1451",
		x"1431", x"11EB", x"0D58", x"06DA", x"FF82", x"F854", x"F277", x"EE55",
		x"EBEE", x"EAE1", x"EACE", x"EB2F", x"EBA2", x"EC0F", x"ECA3", x"EDA0",
		x"EF07", x"F14C", x"F43D", x"F7AC", x"FB11", x"FDDE", x"FF81", x"FFC9",
		x"FEB6", x"FC64", x"F949", x"F613", x"F337", x"F0F7", x"EF8C", x"EF15",
		x"F00A", x"F2E0", x"F7A3", x"FE16", x"054E", x"0C36", x"1135", x"131B",
		x"114C", x"0C68", x"05BE", x"FEAB", x"F80E", x"F252", x"EE0E", x"EBF5",
		x"ECE1", x"F0CA", x"F791", x"002A", x"08A3", x"0F63", x"1357", x"14E4",
		x"14CB", x"1422", x"1389", x"136C", x"13BA", x"144E", x"14DD", x"14E7",
		x"1421", x"12A2", x"1046", x"0D3C", x"09A9", x"05D1", x"0266", x"0000",
		x"FF6A", x"00E9", x"04AF", x"09EE", x"0F5C", x"12EC", x"1317", x"101D",
		x"0B6A", x"0762", x"058D", x"06CC", x"0AA8", x"0F42", x"1263", x"1278",
		x"0EFC", x"08FB", x"01F1", x"FB53", x"F5E2", x"F205", x"EF84", x"EE0E",
		x"ED46", x"ED3F", x"EDFC", x"F061", x"F4BF", x"FB32", x"02F4", x"0A66",
		x"102D", x"138F", x"1497", x"1430", x"139F", x"13A4", x"143E", x"14CF",
		x"147C", x"137E", x"124B", x"11A2", x"11CC", x"12B3", x"13CD", x"1472",
		x"1471", x"141C", x"13BA", x"13EC", x"142E", x"13AF", x"1163", x"0C93",
		x"0579", x"FD87", x"F634", x"F0DC", x"EDE6", x"ECD3", x"ED11", x"EE16",
		x"EFEF", x"F28D", x"F5F0", x"F9C1", x"FD90", x"0107", x"03E4", x"061D",
		x"0829", x"09FA", x"0BC6", x"0D78", x"0F4B", x"112C", x"12E1", x"1444",
		x"1506", x"151C", x"14E2", x"1472", x"1407", x"13EF", x"1436", x"1493",
		x"14D9", x"14B3", x"1419", x"1360", x"12AB", x"1222", x"11D0", x"11F4",
		x"1250", x"1308", x"13D7", x"1487", x"14B1", x"13A3", x"10B1", x"0B21",
		x"0352", x"FAC6", x"F33E", x"EE19", x"EB86", x"EA95", x"EA7C", x"EB0D",
		x"ECAE", x"EFF7", x"F5A0", x"FD36", x"0599", x"0CFD", x"11FB", x"144D",
		x"14C9", x"1487", x"141C", x"13A1", x"12F9", x"1239", x"1124", x"0FB6",
		x"0E2D", x"0C7E", x"0AC9", x"08C5", x"0661", x"0324", x"FEE1", x"F9D1",
		x"F48B", x"F00D", x"ED9D", x"EE0A", x"F189", x"F703", x"FCE0", x"011F",
		x"02B2", x"01AC", x"FEB1", x"FAC3", x"F6DC", x"F38A", x"F148", x"F0E8",
		x"F33C", x"F8B0", x"00A3", x"0909", x"0F78", x"12A4", x"134C", x"12CC",
		x"12CD", x"1314", x"1317", x"115F", x"0CEB", x"05E2", x"FDC2", x"F6DF",
		x"F36A", x"F462", x"F95B", x"00AF", x"0893", x"0EEC", x"12BE", x"13C2",
		x"1287", x"1091", x"0F54", x"0FB2", x"113A", x"130B", x"1497", x"1538",
		x"150D", x"141C", x"12D7", x"1182", x"1050", x"0EF9", x"0D6C", x"0B93",
		x"0939", x"0660", x"032B", x"FFBB", x"FC55", x"F93B", x"F698", x"F496",
		x"F362", x"F2D4", x"F2F9", x"F3E5", x"F531", x"F705", x"F924", x"FBAB",
		x"FEA6", x"0219", x"05E2", x"09B1", x"0D44", x"1027", x"125D", x"13C3",
		x"148C", x"14BF", x"1400", x"1167", x"0C5C", x"0504", x"FCB9", x"F52C",
		x"EF7E", x"EC09", x"EA7F", x"EA4D", x"EB4D", x"EDE4", x"F296", x"F9C3",
		x"0291", x"0B1A", x"116B", x"149B", x"153A", x"14C8", x"1461", x"1420",
		x"13CA", x"12DE", x"1105", x"0DE1", x"0907", x"0275", x"FB1A", x"F412",
		x"EEDA", x"EC4C", x"EC68", x"EEB5", x"F25D", x"F6A1", x"FAE1", x"FEB7",
		x"01E6", x"045C", x"061C", x"06CF", x"0650", x"047E", x"0147", x"FD40",
		x"F922", x"F580", x"F31F", x"F282", x"F44E", x"F8BF", x"FF73", x"0701"
	);

	constant q_vals : vals := (
		x"EB93", x"ECD7", x"EEF9", x"F227", x"F67B", x"FBE9", x"0203", x"0835",
		x"0DCB", x"11EC", x"13C2", x"12B6", x"0E85", x"07CA", x"FFD8", x"F829",
		x"F1DE", x"EDAD", x"EBAC", x"EC03", x"EF10", x"F4C8", x"FC78", x"04F1",
		x"0C8C", x"11A7", x"1397", x"1290", x"0FE6", x"0D38", x"0BD2", x"0C1D",
		x"0DB3", x"0FD5", x"11EF", x"1399", x"149F", x"1503", x"14AD", x"1361",
		x"1080", x"0BA4", x"04E0", x"FCEB", x"F527", x"EF0D", x"EC55", x"EDCF",
		x"F39C", x"FBE5", x"0499", x"0BEC", x"1108", x"140A", x"153E", x"14ED",
		x"1328", x"0FE7", x"0AB4", x"0371", x"FB4B", x"F3A7", x"EE48", x"EBC5",
		x"EBCD", x"ED28", x"EED5", x"F05A", x"F15B", x"F1F6", x"F245", x"F25A",
		x"F241", x"F233", x"F1E9", x"F114", x"EF90", x"EDB0", x"EBF1", x"EB53",
		x"ECAA", x"F035", x"F5F1", x"FD66", x"051E", x"0BC9", x"10A2", x"1391",
		x"14F8", x"1552", x"1548", x"14FE", x"1496", x"13A0", x"11CF", x"0EA0",
		x"0A01", x"039B", x"FC3A", x"F4DE", x"EF4C", x"EC96", x"ECBA", x"EEEC",
		x"F16D", x"F31E", x"F32B", x"F1E0", x"EFD7", x"EDBF", x"EC12", x"EB01",
		x"EA6B", x"EAB6", x"EC73", x"F053", x"F678", x"FE3A", x"0659", x"0D44",
		x"1220", x"1488", x"1538", x"1520", x"14DE", x"1490", x"13C8", x"1246",
		x"0F85", x"0B85", x"05DD", x"FF17", x"F7FC", x"F1E9", x"EDC6", x"EC31",
		x"ED17", x"F011", x"F43F", x"F8D9", x"FD11", x"0049", x"0273", x"03E3",
		x"053D", x"06D4", x"08CB", x"0AF1", x"0D44", x"0F7E", x"116B", x"12C4",
		x"13D2", x"1460", x"14BA", x"14DC", x"14D2", x"14BD", x"1428", x"134A",
		x"11C5", x"0FB9", x"0CDB", x"08F1", x"03A8", x"FD4F", x"F689", x"F093",
		x"ECCD", x"EC02", x"EE89", x"F3C2", x"FAC6", x"0254", x"095D", x"0F00",
		x"12C4", x"1443", x"1310", x"0EF1", x"081B", x"FF84", x"F6C0", x"EFE0",
		x"EC2E", x"EBC2", x"ED57", x"EF2E", x"EFDB", x"EF20", x"ED79", x"EC46",
		x"ECFC", x"F083", x"F6F7", x"FF7B", x"084D", x"0F3B", x"129B", x"11BB",
		x"0D19", x"0678", x"FFAB", x"FA77", x"F814", x"F952", x"FDE6", x"049B",
		x"0B73", x"105E", x"1291", x"125D", x"10D6", x"0FA1", x"0FDC", x"116F",
		x"12DD", x"11C1", x"0CF9", x"053B", x"FCB7", x"F58E", x"F09D", x"EDDA",
		x"ECA6", x"EC60", x"EC44", x"EBCB", x"EB49", x"EB42", x"EC94", x"EFF4",
		x"F585", x"FCCB", x"04B1", x"0BE3", x"1149", x"1461", x"1533", x"145E",
		x"12B6", x"10CF", x"0F2C", x"0D82", x"0BD9", x"0A1F", x"085A", x"06BB",
		x"0508", x"039F", x"0219", x"0021", x"FD50", x"F988", x"F515", x"F0A0",
		x"ED73", x"ECC0", x"EF2C", x"F466", x"FB24", x"0196", x"0632", x"0807",
		x"0687", x"026C", x"FC7E", x"F615", x"F09D", x"EDC3", x"EEA5", x"F370",
		x"FAB9", x"02A3", x"0983", x"0ED4", x"126E", x"143B", x"13AD", x"0FFE",
		x"095C", x"008A", x"F776", x"F031", x"EC32", x"EB93", x"ECFE", x"EEA6",
		x"EF0A", x"EE01", x"ECAB", x"ECC9", x"EFAC", x"F5B6", x"FD92", x"04F6",
		x"0A2D", x"0C8B", x"0C5F", x"0A07", x"0625", x"019D", x"FD5A", x"FA90",
		x"F9EC", x"FBB7", x"FFCC", x"0591", x"0BB5", x"109C", x"12F2", x"118F",
		x"0CE5", x"05CD", x"FDC3", x"F62F", x"F03E", x"EC9B", x"EB8E", x"ED3F",
		x"F0F1", x"F5CB", x"FAB2", x"FEEB", x"0226", x"0497", x"066C", x"0830",
		x"09FA", x"0BDF", x"0DF5", x"1019", x"1232", x"1404", x"1516", x"1568",
		x"1566", x"1536", x"1510", x"14DA", x"14B0", x"14A4", x"14B2", x"1473",
		x"1380", x"1173", x"0DA7", x"07AC", x"FFDC", x"F782", x"F0B0", x"ECEF",
		x"EC4E", x"ED4F", x"EE22", x"EE0E", x"ED52", x"ED2E", x"EF0A", x"F3D6",
		x"FB0E", x"02E5", x"0900", x"0B50", x"0937", x"036A", x"FBC5", x"F475",
		x"EF10", x"EC91", x"ECDE", x"EEBF", x"F0FA", x"F237", x"F1E3", x"F045",
		x"EE2C", x"EC87", x"EBA1", x"EBD9", x"EDD4", x"F1FB", x"F87B", x"009F",
		x"089F", x"0F11", x"132F", x"150E", x"1577", x"153F", x"14F7", x"14BB",
		x"1448", x"1368", x"11E8", x"1057", x"0F38", x"0EFC", x"0F8A", x"10B2",
		x"1212", x"1367", x"146F", x"1505", x"14C8", x"13E6", x"125E", x"1048",
		x"0DD2", x"0B36", x"08F0", x"0794", x"07B1", x"096B", x"0C62", x"0FD4",
		x"1250", x"12A1", x"0FE3", x"0A71", x"038A", x"FCAA", x"F713", x"F324",
		x"F0CB", x"EF67", x"EE90", x"EDD6", x"ED0D", x"EC2E", x"EB67", x"EB0A",
		x"EB50", x"EC68", x"EDF9", x"EF59", x"F001", x"EFA0", x"EE89", x"ED0B",
		x"EBF9", x"ECAE", x"EFDB", x"F596", x"FD1D", x"04E2", x"0B86", x"1061",
		x"1333", x"1460", x"1492", x"144E", x"140E", x"1420", x"147B", x"14AB",
		x"1402", x"11ED", x"0DA0", x"0747", x"FF83", x"F78A", x"F0F5", x"ED1E",
		x"ECDF", x"F07E", x"F70A", x"FF0F", x"06C8", x"0CDF", x"10E2", x"12F3",
		x"13A1", x"1318", x"117C", x"0F0C", x"0C28", x"0962", x"0781", x"0713",
		x"089C", x"0BC3", x"0FB4", x"1291", x"1299", x"0EFF", x"08A4", x"016C",
		x"FB10", x"F68A", x"F3D5", x"F253", x"F170", x"F095", x"EF1E", x"ED52",
		x"EBC0", x"EB9E", x"EDBA", x"F290", x"F96E", x"0161", x"08BD", x"0E95",
		x"1238", x"13CB", x"13C6", x"12C3", x"1126", x"0EFD", x"0C7B", x"09CA",
		x"075F", x"05D6", x"0557", x"0626", x"07DC", x"0A46", x"0CD2", x"0F7E",
		x"11EB", x"13A9", x"145D", x"1359", x"104F", x"0B1C", x"0433", x"FC56",
		x"F4C1", x"EEED", x"EBF6", x"EC54", x"EFED", x"F600", x"FD7F", x"04FC",
		x"0B5A", x"1004", x"12EB", x"146C", x"14D0", x"147A", x"13E5", x"1355",
		x"12EE", x"1243", x"110D", x"0EF8", x"0C13", x"0864", x"041C", x"FFFF",
		x"FCCA", x"FB82", x"FCA0", x"0047", x"060F", x"0C6A", x"114D", x"12AD",
		x"107C", x"0C48", x"08D0", x"07EE", x"0A2B", x"0E4C", x"11D5", x"128A",
		x"0F6B", x"09B0", x"03DF", x"00C7", x"01BD", x"063E", x"0C16", x"10B6",
		x"1211", x"0FD3", x"0B94", x"0811", x"0732", x"099E", x"0DE4", x"115D",
		x"11F0", x"0EC3", x"090B", x"0308", x"FEC6", x"FD0A", x"FDF5", x"00C2",
		x"04A9", x"08C8", x"0C5E", x"0EAA", x"0FC2", x"0FBB", x"0EB2", x"0CB3",
		x"09D4", x"069E", x"0378", x"0100", x"FF58", x"FECD", x"FF58", x"00DE",
		x"0346", x"0637", x"0961", x"0C60", x"0F1C", x"1122", x"129E", x"13A7",
		x"1463", x"14C6", x"1503", x"14FD", x"148C", x"13C1", x"1236", x"1007",
		x"0D93", x"0AD0", x"081C", x"05E1", x"0456", x"03BD", x"0441", x"05A4",
		x"07B7", x"0A5D", x"0D14", x"0F79", x"1125", x"1216", x"128C", x"128B",
		x"1254", x"1162", x"0FC0", x"0D63", x"0A1B", x"05F7", x"00D0", x"FB1B",
		x"F53C", x"F062", x"ED10", x"EC15", x"EDD1", x"F26D", x"F96D", x"01B9",
		x"09C5", x"0FFC", x"1376", x"13D9", x"1172", x"0D13", x"07B7", x"024E",
		x"FD83", x"F9C8", x"F6D0", x"F47E", x"F28E", x"F0DC", x"EF97", x"EE5D",
		x"ED7D", x"ECB6", x"EC20", x"EBC5", x"EB66", x"EB27", x"EB28", x"EC48",
		x"EF94", x"F599", x"FDE7", x"06BB", x"0DE8", x"1250", x"1446", x"14DB",
		x"14DC", x"1486", x"12E5", x"0F4F", x"094E", x"015B", x"F8CA", x"F1B1",
		x"EE18", x"EF12", x"F463", x"FC7A", x"0523", x"0C5E", x"115F", x"142D",
		x"1532", x"1515", x"141B", x"11A9", x"0D18", x"0655", x"FDE1", x"F5E3",
		x"F04C", x"EE90", x"F0B9", x"F640", x"FDFD", x"0617", x"0D23", x"11F1",
		x"1425", x"1448", x"137A", x"12F3", x"133F", x"141D", x"14D1", x"14AD",
		x"13FA", x"133D", x"12F8", x"1336", x"13CF", x"1475", x"14E2", x"14E0",
		x"1449", x"132B", x"11B6", x"101B", x"0E73", x"0CDD", x"0B05", x"08BF",
		x"064A", x"0376", x"006E", x"FD78", x"FA82", x"F7D2", x"F59C", x"F396",
		x"F1F4", x"F06C", x"EEFC", x"ED6D", x"EC2F", x"EB54", x"EB25", x"EB7E",
		x"EC15", x"ECA1", x"ED0B", x"ED15", x"EC9C", x"EBEE", x"EB4D", x"EB0D",
		x"EB5B", x"EBEB", x"EC4B", x"EC10", x"EB90", x"EB86", x"ED07", x"F0D3",
		x"F71D", x"FF36", x"078A", x"0E85", x"12F7", x"142A", x"1257", x"0E0F",
		x"07E9", x"00A8", x"F93A", x"F2B0", x"EE17", x"EC3B", x"ED55", x"F12A",
		x"F744", x"FEB3", x"060A", x"0C53", x"10BA", x"1364", x"14AF", x"1524",
		x"153C", x"14F2", x"148C", x"13F0", x"12FB", x"115E", x"0EE1", x"0B65",
		x"0745", x"0325", x"FFD8", x"FE25", x"FEA1", x"019D", x"069F", x"0C80",
		x"1158", x"136A", x"1200", x"0E35", x"09E8", x"072A", x"06F4", x"096F",
		x"0D6F", x"115C", x"1336", x"117F", x"0BF9", x"03A1", x"FA51", x"F24A",
		x"ED6F", x"EC8B", x"EF09", x"F383", x"F850", x"FBA1", x"FC6D", x"FA4C",
		x"F5EF", x"F0EA", x"ED9B", x"ED73", x"F09B", x"F59E", x"FA53", x"FD43",
		x"FD9F", x"FB94", x"F7E2", x"F3B8", x"F008", x"ED78", x"EC22", x"EC46",
		x"EDC0", x"F068", x"F396", x"F6EE", x"F9E0", x"FBE7", x"FC4C", x"FA86",
		x"F6CD", x"F214", x"EE21", x"EC99", x"EE3D", x"F2AB", x"F8BA", x"FF19",
		x"04B4", x"0921", x"0C31", x"0E19", x"0F60", x"104D", x"114E", x"1244",
		x"133C", x"13F8", x"1473", x"14AC", x"1422", x"1347", x"1241", x"119C",
		x"1175", x"11D7", x"12D6", x"13D5", x"14AA", x"14F8", x"14BA", x"1465",
		x"1439", x"1464", x"14A9", x"14D7", x"1491", x"13C0", x"12DE", x"1257",
		x"1294", x"136F", x"1443", x"1463", x"12B4", x"0E88", x"07D1", x"FF6C",
		x"F6F7", x"F04B", x"ECD7", x"ED0E", x"F097", x"F662", x"FD12", x"03A6",
		x"08FD", x"0CC2", x"0EC1", x"0F61", x"0E7E", x"0C86", x"098D", x"05DD",
		x"01D4", x"FDB2", x"F9EF", x"F6DF", x"F497", x"F2ED", x"F1A7", x"F060",
		x"EF07", x"ED74", x"EC06", x"EAFB", x"EAAA", x"EB3B", x"EC58", x"EDCA",
		x"EEDD", x"EF31", x"EE4F", x"ECF2", x"EC2C", x"ED5B", x"F139", x"F7D9",
		x"FFEA", x"0786", x"0D05", x"0F8C", x"0F52", x"0D04", x"094F", x"04C3",
		x"0054", x"FD17", x"FC0E", x"FDFF", x"029E", x"0902", x"0F12", x"1286",
		x"125A", x"0F5D", x"0B9F", x"0958", x"09A7", x"0C61", x"0FF4", x"126A",
		x"121C", x"0E9A", x"087C", x"0158", x"FAA5", x"F53C", x"F17C", x"EF37",
		x"EDF7", x"ED3D", x"ECA6", x"EC3C", x"EC1F", x"EC87", x"ED44", x"EE5B",
		x"EFE5", x"F1E8", x"F492", x"F7AB", x"FB10", x"FE48", x"0139", x"0393",
		x"0590", x"0754", x"093A", x"0B6D", x"0DCD", x"1047", x"127E", x"1424",
		x"1507", x"153D", x"1533", x"1529", x"154A", x"1544", x"144B", x"1158",
		x"0C00", x"04BC", x"FCB0", x"F552", x"EFDC", x"ECA5", x"EB99", x"EC1F",
		x"EDAE", x"EFD3", x"F28F", x"F564", x"F78A", x"F82C", x"F6EE", x"F3F2",
		x"F046", x"ED6B", x"ED0B", x"EFE5", x"F5F4", x"FDCA", x"05FC", x"0D0D",
		x"11DA", x"13BC", x"12B7", x"0F2C", x"09EA", x"03C5", x"FD93", x"F7EC",
		x"F364", x"F036", x"EE32", x"ED1F", x"EC90", x"EC45", x"EBFE", x"EBF0",
		x"EC1C", x"ECC0", x"EDF5", x"EFB2", x"F21E", x"F4EC", x"F7F0", x"FAD9",
		x"FD75", x"FF95", x"014A", x"02BE", x"0460", x"0695", x"09E6", x"0DD3",
		x"114E", x"12EE", x"11B3", x"0D68", x"06A5", x"FF0A", x"F87A", x"F4D2",
		x"F50F", x"F91D", x"FFB6", x"073D", x"0DC9", x"11E3", x"131C", x"1213",
		x"1053", x"0F6A", x"0FF1", x"11CB", x"13B5", x"14D0", x"1533", x"1532",
		x"154B", x"14F3", x"13A1", x"106F", x"0B24", x"03B7", x"FB66", x"F380",
		x"EE10", x"EC1E", x"EE08", x"F32E", x"FA8D", x"0271", x"09AA", x"0F2B",
		x"1299", x"142D", x"1474", x"13D4", x"1293", x"10AC", x"0E21", x"0B6C",
		x"08FC", x"079C", x"079E", x"08DC", x"0B13", x"0DBF", x"1058", x"1276",
		x"13FC", x"14D4", x"14F9", x"14C2", x"143A", x"1399", x"12A7", x"110D",
		x"0E6C", x"0A76", x"04E7", x"FE18", x"F6FC", x"F0D1", x"ED25", x"EC8C",
		x"EE93", x"F20C", x"F560", x"F74F", x"F749", x"F573", x"F29F", x"EFB5",
		x"ED3F", x"EB9B", x"EACE", x"EAC4", x"EB71", x"EC9F", x"EE05", x"EFAA",
		x"F1B5", x"F3DA", x"F585", x"F658", x"F659", x"F5CC", x"F4CE", x"F378",
		x"F1B0", x"EF88", x"ED80", x"EC56", x"ECBE", x"EFA3", x"F501", x"FC30",
		x"03E3", x"0ADC", x"101C", x"1327", x"1498", x"14F9", x"14D1", x"140E",
		x"129E", x"106F", x"0DA2", x"0A79", x"0713", x"0397", x"002C", x"FD23",
		x"FA66", x"F85C", x"F6C0", x"F5A6", x"F505", x"F4E3", x"F532", x"F5E2",
		x"F70C", x"F900", x"FC0C", x"00AF", x"0660", x"0C2A", x"10DB", x"1342",
		x"12E0", x"0FB1", x"0AB4", x"04FC", x"FF85", x"FB3C", x"F879", x"F770",
		x"F7BE", x"F993", x"FC83", x"00DF", x"065B", x"0BE7", x"10B3", x"1362",
		x"133B", x"105F", x"0B2E", x"04C5", x"FE8C", x"F954", x"F5AB", x"F3D7",
		x"F396", x"F487", x"F6BE", x"FA5C", x"FFBD", x"064D", x"0C22", x"0E92",
		x"0C8C", x"07F4", x"04D1", x"05DA", x"0AC9", x"10B5", x"14D3", x"1625",
		x"15D8", x"1522", x"14A0", x"13B7", x"11E3", x"0EB9", x"09E5", x"03C4",
		x"FCE3", x"F615", x"F079", x"ECFC", x"EC1A", x"EDB9", x"F15F", x"F5DA",
		x"FA59", x"FDEB", x"0062", x"01FA", x"0365", x"0522", x"07B6", x"0B29",
		x"0EDB", x"121B", x"1393", x"1237", x"0DDA", x"0726", x"FF7A", x"F86B",
		x"F348", x"F013", x"EE73", x"ED83", x"ECBB", x"EBEF", x"EB28", x"EAE3",
		x"EB45", x"ED1F", x"F0B2", x"F643", x"FDA0", x"0592", x"0CB8", x"11B0",
		x"13A2", x"1275", x"0EA5", x"08F1", x"01F7", x"FA87", x"F3BF", x"EE9D",
		x"EBE3", x"EC0C", x"EEFB", x"F42C", x"FAEE", x"0259", x"0968", x"0F2D",
		x"12E7", x"141C", x"126E", x"0E21", x"07DA", x"007C", x"F904", x"F276",
		x"EDAF", x"EB85", x"EC5E", x"F006", x"F59B", x"FC77", x"0392", x"0A2F",
		x"0F87", x"12B2", x"12A9", x"0EF4", x"0848", x"000A", x"F828", x"F1DB",
		x"EDAA", x"EB5E", x"EABA", x"EBB8", x"EE53", x"F2DE", x"F975", x"01C1",
		x"0A2C", x"108C", x"1364", x"1256", x"0E43", x"0872", x"018E", x"FA5C",
		x"F3CF", x"EF05", x"EC9F", x"ECD4", x"EF83", x"F460", x"FAC7", x"0225",
		x"0931", x"0EF0", x"1282", x"1374", x"11AF", x"0DAF", x"07FA", x"011C",
		x"FA1B", x"F3BB", x"EEB1", x"EC41", x"ED52", x"F268", x"FAA5", x"03DA",
		x"0BBA", x"111C", x"1445", x"1577", x"14EB", x"122D", x"0D28", x"0647",
		x"FE64", x"F6A0", x"F02C", x"EBEA", x"EA04", x"EA96", x"ED5E", x"F266",
		x"F9B0", x"024F", x"0AA3", x"10DA", x"137A", x"125D", x"0E1B", x"0816",
		x"010E", x"FA0D", x"F3C2", x"EED5", x"EC32", x"EC9E", x"F020", x"F65A",
		x"FE29", x"0609", x"0C94", x"113A", x"13F3", x"1523", x"14EC", x"13A9",
		x"11D4", x"0FBC", x"0DDC", x"0C51", x"0AED", x"096A", x"07C4", x"05FC",
		x"03EB", x"01AC", x"FF0B", x"FBFF", x"F87D", x"F4AA", x"F0DE", x"EDAF",
		x"EBF6", x"EC73", x"EF8D", x"F522", x"FC86", x"048F", x"0BEF", x"114B",
		x"13BA", x"135D", x"107D", x"0BD6", x"058B", x"FE48", x"F6E7", x"F0C8",
		x"ED7D", x"EDFB", x"F233", x"F8DC", x"FFE8", x"05BA", x"08BC", x"082C",
		x"03B3", x"FC7A", x"F4E2", x"EF55", x"ED1A", x"ED8B", x"EEF7", x"EF96",
		x"EEED", x"EDB4", x"EDC0", x"F0BA", x"F6EE", x"FEE1", x"0605", x"09B5",
		x"088B", x"02FA", x"FB02", x"F363", x"EE73", x"ECBB", x"ED73", x"EED4",
		x"EF4E", x"EE8B", x"ED40", x"ECFB", x"EF7C", x"F561", x"FD77", x"05AF",
		x"0C3A", x"1069", x"12C9", x"140F", x"14B8", x"1510", x"152E", x"1543",
		x"151C", x"1495", x"13C6", x"128D", x"10E7", x"0EFA", x"0CF8", x"0AEB",
		x"08F8", x"06DE", x"0481", x"01FD", x"FF4D", x"FCB9", x"FA01", x"F73D",
		x"F4A9", x"F246", x"F080", x"EF2F", x"EE3A", x"ED86", x"ECCE", x"EBD5",
		x"EAFF", x"EB5E", x"EDEB", x"F391", x"FBBA", x"0481", x"0C12", x"1154",
		x"142F", x"1572", x"153C", x"134C", x"0F44", x"090A", x"0162", x"F961",
		x"F285", x"EDE7", x"EBF4", x"EC8D", x"EF9D", x"F4D9", x"FC2F", x"0489",
		x"0C68", x"11BE", x"1355", x"1115", x"0C1E", x"05A9", x"FEAF", x"F7F4",
		x"F21E", x"EDE5", x"EC25", x"ED9B", x"F29B", x"FA46", x"02C1", x"0A4A",
		x"0FC9", x"12F9", x"1468", x"14E5", x"150D", x"1540", x"1562", x"1503",
		x"13F3", x"127A", x"10D6", x"0F5D", x"0E93", x"0E80", x"0F1E", x"105D",
		x"11DE", x"134F", x"1437", x"1412", x"1263", x"0F10", x"0A23", x"039C",
		x"FC2E", x"F512", x"EF9E", x"ECEA", x"ED88", x"F142", x"F75E", x"FECB",
		x"0679", x"0CFE", x"11A2", x"140C", x"1478", x"1383", x"11A5", x"0F49",
		x"0C9A", x"0A1B", x"0821", x"0702", x"06FE", x"0829", x"0A31", x"0CED",
		x"0FBD", x"1224", x"13C2", x"14BA", x"14F4", x"13FF", x"1098", x"0A5E",
		x"020E", x"F9A4", x"F2C6", x"EDF7", x"EB27", x"E9E0", x"EA50", x"ECBD",
		x"F168", x"F814", x"0034", x"089B", x"0FA0", x"13B5", x"1423", x"110D",
		x"0B3E", x"03A2", x"FB52", x"F396", x"EDE3", x"EB04", x"EA45", x"EA96",
		x"EAF1", x"EB16", x"EBA3", x"ECC9", x"EE54", x"EFA1", x"F04A", x"F013",
		x"EF2A", x"EDD5", x"EC84", x"EB70", x"EAE5", x"EABA", x"EAD5", x"EAE0",
		x"EAEE", x"EB02", x"EB47", x"EBFC", x"ED1A", x"EEA0", x"EFC4", x"F052",
		x"F008", x"EF14", x"EDAC", x"EC63", x"EB50", x"EAA1", x"EA74", x"EAFB",
		x"EC18", x"EDDA", x"F005", x"F24E", x"F473", x"F698", x"F842", x"F915",
		x"F900", x"F7CD", x"F5C7", x"F33C", x"F0ED", x"EF14", x"ED82", x"EC59",
		x"EB9A", x"EB84", x"EC24", x"ED79", x"EF65", x"F1F5", x"F50A", x"F83D",
		x"FB42", x"FDC6", x"FFDA", x"017C", x"02DE", x"0460", x"06AF", x"0A0D",
		x"0DD2", x"1104", x"12E8", x"12A9", x"0FFB", x"0AE7", x"040F", x"FCC2",
		x"F647", x"F16E", x"EE2D", x"EC3C", x"EB43", x"EABE", x"EAD7", x"EB2D",
		x"EBAB", x"EC0A", x"EC75", x"ECF4", x"EDCA", x"EEFA", x"F0D2", x"F349",
		x"F6BC", x"FB01", x"0018", x"058B", x"0B3C", x"102D", x"1364", x"13E0",
		x"110B", x"0B4D", x"0354", x"FABA", x"F315", x"EE17", x"EC89", x"EE1E",
		x"F154", x"F4AF", x"F656", x"F5BE", x"F2FE", x"EF70", x"ECC0", x"EC7B",
		x"EF94", x"F5E1", x"FE6B", x"0747", x"0E64", x"1234", x"1252", x"0F16",
		x"09CD", x"046C", x"00DC", x"009C", x"03EE", x"097B", x"0F32", x"12C1",
		x"12CE", x"0FD0", x"0B98", x"089D", x"0881", x"0B58", x"0F89", x"128B",
		x"123F", x"0E3F", x"080F", x"01E5", x"FD5D", x"FB3E", x"FB55", x"FD59",
		x"00D3", x"0500", x"097C", x"0DD1", x"1178", x"13A6", x"13C9", x"118A",
		x"0C9C", x"05DB", x"FE40", x"F719", x"F1A9", x"EE35", x"EC42", x"EB40",
		x"EABF", x"EAB2", x"EAD9", x"EB33", x"EBB6", x"EC77", x"ED7F", x"EEE1",
		x"F07D", x"F24D", x"F45B", x"F6C5", x"F9A5", x"FD02", x"00BB", x"045D",
		x"07AE", x"0A9D", x"0D10", x"0EF2", x"0FA1", x"0EC3", x"0C24", x"07B2",
		x"01D4", x"FB0E", x"F42D", x"EEFC", x"ECBC", x"EE07", x"F2A8", x"F94E",
		x"00AA", x"079F", x"0D76", x"11C1", x"1400", x"137C", x"0FAE", x"08DE",
		x"0004", x"F6FE", x"EFDB", x"EBF4", x"EAC3", x"EB3B", x"EBC0", x"EBB7",
		x"EBA6", x"EC8B", x"EF7E", x"F4D6", x"FC54", x"047C", x"0BCD", x"1125",
		x"141E", x"1506", x"14A9", x"1398", x"12C0", x"12A0", x"135E", x"1447",
		x"13FE", x"11B1", x"0D02", x"067B", x"FF06", x"F7CC", x"F210", x"EEF5",
		x"EEE6", x"F219", x"F80F", x"FFA7", x"07C9", x"0EB2", x"1309", x"13EF",
		x"125D", x"0FB5", x"0D86", x"0C50", x"0BAF", x"0AD4", x"08EA", x"05A5",
		x"0081", x"F9FC", x"F37A", x"EEAE", x"ECD0", x"EE41", x"F1F4", x"F66E",
		x"FA38", x"FC5D", x"FCB9", x"FB9A", x"F97A", x"F6B5", x"F3AA", x"F0C2",
		x"EE3F", x"EC60", x"EB4C", x"EB1C", x"EBBF", x"ECE8", x"EE0C", x"EE7B",
		x"EDF8", x"ECCB", x"EC36", x"ED4D", x"F0D1", x"F68F", x"FDD7", x"056B",
		x"0B9B", x"0F1D", x"0EFA", x"0B1C", x"049C", x"FCBF", x"F533", x"EF66",
		x"EC88", x"EC79", x"EEA9", x"F1C1", x"F450", x"F5D9", x"F6B1", x"F7E2",
		x"FA03", x"FDA0", x"028F", x"0883", x"0E3C", x"1256", x"1373", x"1156",
		x"0CCC", x"0781", x"0342", x"011C", x"0125", x"033A", x"066E", x"0A11",
		x"0D41", x"0FAE", x"10F7", x"1117", x"0FD7", x"0D69", x"0A28", x"0658",
		x"02BB", x"0050", x"FFFD", x"024D", x"06DA", x"0C7D", x"1139", x"12FB",
		x"110D", x"0C5E", x"0776", x"04A1", x"0547", x"08E4", x"0DBF", x"11B0",
		x"12EB", x"109B", x"0B81", x"04E4", x"FE9D", x"F98C", x"F614", x"F3EF",
		x"F285", x"F163", x"F02F", x"EF13", x"EDE1", x"EC9A", x"EB9B", x"EB19",
		x"EB26", x"EBA3", x"EC47", x"ECA0", x"ECC4", x"EC89", x"EC16", x"EBA3",
		x"EB77", x"EBD5", x"EC89", x"ED2B", x"ED4D", x"ECF9", x"EC36", x"EB6D",
		x"EB29", x"EB8D", x"EC73", x"ED01", x"ECA7", x"EBDC", x"EBD2", x"EDE6",
		x"F273", x"F934", x"010C", x"089B", x"0E7D", x"1127", x"102E", x"0B97",
		x"048D", x"FC81", x"F4F3", x"EF5E", x"EC41", x"EBB0", x"EC6D", x"ED2E",
		x"ED1A", x"EC40", x"EB4E", x"EAF0", x"EB8E", x"ECEC", x"EEA8", x"F0AE",
		x"F2DB", x"F4FA", x"F703", x"F932", x"FB91", x"FE28", x"00CC", x"03A4",
		x"06AC", x"09C4", x"0C87", x"0EC3", x"1067", x"1189", x"1211", x"11EA",
		x"110E", x"0F78", x"0D26", x"0A3C", x"0728", x"0484", x"02EB", x"0293",
		x"03C3", x"0679", x"09F1", x"0D7E", x"1049", x"1235", x"133D", x"12AD",
		x"0FA5", x"09AD", x"01B9", x"F963", x"F283", x"EDF2", x"EB6C", x"EAA2",
		x"EABA", x"EB7B", x"ED3D", x"F0DB", x"F6BE", x"FEA3", x"06FA", x"0DDB",
		x"1255", x"146D", x"1505", x"14EA", x"1492", x"1408", x"1351", x"127B",
		x"116E", x"0FEC", x"0E24", x"0BDD", x"0973", x"06EF", x"0463", x"01DB",
		x"FF2E", x"FC68", x"F9A6", x"F6CB", x"F3F6", x"F130", x"EF0D", x"ED7F",
		x"ECC4", x"ECF5", x"EDC7", x"EF9B", x"F254", x"F5F3", x"F971", x"FC2E",
		x"FD2E", x"FBD5", x"F848", x"F385", x"EF3A", x"ED8B", x"EF83", x"F4AA",
		x"FA6C", x"FE47", x"FE6C", x"FAC8", x"F510", x"EFC0", x"ED3B", x"EE5E",
		x"F23A", x"F65A", x"F891", x"F7C5", x"F455", x"F027", x"ED75", x"EE0D",
		x"F257", x"F8FC", x"FFF1", x"05D6", x"0A3D", x"0D10", x"0EB3", x"0F8F",
		x"104E", x"113E", x"1281", x"13D1", x"14CC", x"1532", x"14F2", x"1417",
		x"12F6", x"11EE", x"1170", x"1193", x"124D", x"1311", x"13F0", x"1491",
		x"14FE", x"152D", x"151F", x"14F2", x"14BC", x"14A3", x"14C6", x"14FC",
		x"1530", x"14D6", x"13AA", x"10E0", x"0C06", x"0514", x"FCBE", x"F4FF",
		x"EF3D", x"EC69", x"EBF3", x"EC59", x"EC8B", x"EC41", x"EC29", x"EDA6",
		x"F19F", x"F83D", x"003B", x"07DA", x"0D52", x"1014", x"10B1", x"0FAA",
		x"0D28", x"0987", x"0526", x"0090", x"FC77", x"F95F", x"F73D", x"F5C7",
		x"F4C7", x"F3B2", x"F24D", x"F02D", x"EDC9", x"EBF2", x"EC04", x"EEBE",
		x"F436", x"FB66", x"031C", x"0A2E", x"0F63", x"1280", x"13CE", x"13BE",
		x"12C6", x"10E0", x"0E04", x"0A9D", x"0793", x"05AA", x"0583", x"0724",
		x"09E7", x"0D11", x"1001", x"128C", x"1471", x"1522", x"13DD", x"0FDC",
		x"092E", x"00D1", x"F86E", x"F1B2", x"ED5A", x"EB36", x"EA86", x"EACF",
		x"EC81", x"F02A", x"F5D7", x"FD68", x"0571", x"0C94", x"1176", x"13E8",
		x"1488", x"1443", x"135B", x"11AB", x"0F0C", x"0BB9", x"07F6", x"0459",
		x"00F7", x"FDE1", x"FAF0", x"F842", x"F5D6", x"F3F1", x"F2B6", x"F220",
		x"F286", x"F3BD", x"F5BA", x"F89B", x"FBF4", x"FF4F", x"0206", x"03AB",
		x"03FB", x"02EB", x"00A4", x"FD57", x"F98F", x"F623", x"F376", x"F21F",
		x"F1FD", x"F32A", x"F588", x"F8E3", x"FCD8", x"0090", x"036E", x"0463",
		x"0303", x"FF41", x"F996", x"F36B", x"EEBB", x"ECC1", x"EDD7", x"F132",
		x"F52E", x"F858", x"F9D1", x"F94B", x"F733", x"F448", x"F13C", x"EE80",
		x"EC69", x"EB2F", x"EAD8", x"EB20", x"EBC7", x"EC61", x"ECF4", x"EDBF",
		x"EF09", x"F106", x"F382", x"F5F9", x"F84F", x"FA57", x"FC78", x"FED8",
		x"018C", x"0482", x"077F", x"0A34", x"0CB0", x"0EF5", x"1103", x"12B8",
		x"13E6", x"145B", x"145C", x"143B", x"1416", x"13C4", x"1341", x"1215",
		x"0FBE", x"0BDC", x"0660", x"FFA1", x"F82B", x"F1AA", x"ED74", x"EC6D",
		x"EE2B", x"F110", x"F369", x"F41E", x"F2F2", x"F059", x"EDFC", x"ED9A",
		x"F092", x"F6C5", x"FEF8", x"0760", x"0E73", x"12C5", x"13EA", x"11E3",
		x"0D86", x"07E3", x"01C4", x"FC07", x"F73E", x"F394", x"F13A", x"EFF3",
		x"EF20", x"EE3C", x"ED17", x"EBF6", x"EBCB", x"EDA8", x"F241", x"F921",
		x"014D", x"0947", x"0F7C", x"1353", x"14B5", x"147A", x"1368", x"11C0",
		x"0FB6", x"0D37", x"0AEE", x"09AF", x"0A26", x"0C49", x"0F89", x"12B9",
		x"142E", x"12E0", x"0E67", x"0712", x"FE31", x"F5A7", x"EF8D", x"ED14",
		x"EE98", x"F2F1", x"F8C8", x"FE56", x"0222", x"0304", x"0082", x"FB78",
		x"F559", x"F015", x"ED20", x"ED80", x"F0A0", x"F5B8", x"FB3D", x"FFF1",
		x"0362", x"05AE", x"075E", x"08DF", x"0A6C", x"0BEB", x"0D58", x"0EB2",
		x"0FEC", x"1126", x"1266", x"1372", x"1473", x"1504", x"1436", x"1147",
		x"0BCC", x"0453", x"FC55", x"F51C", x"EFAA", x"EC4A", x"EACD", x"EA84",
		x"EABA", x"EADA", x"EAA1", x"EA9A", x"EB86", x"EDD1", x"F1DF", x"F7A5",
		x"FF0D", x"071C", x"0E04", x"122F", x"12E6", x"11A4", x"1029", x"1001",
		x"1101", x"125E", x"1250", x"0F6F", x"098D", x"01E4", x"FAE8", x"F6FC",
		x"F780", x"FC38", x"037E", x"0B2F", x"10E3", x"1385", x"1324", x"10C2",
		x"0DEB", x"0BD1", x"0B57", x"0CAE", x"0F00", x"11B7", x"13C9", x"14B8",
		x"13FA", x"1134", x"0CA0", x"066C", x"FF5F", x"F845", x"F21F", x"EDE9",
		x"EBF7", x"EBF2", x"ED38", x"EF21", x"F124", x"F2AF", x"F3BB", x"F441",
		x"F457", x"F402", x"F366", x"F259", x"F11E", x"EFD5", x"EE5A", x"ED02",
		x"EC01", x"EB83", x"EBC0", x"ECD3", x"EE65", x"F052", x"F1E2", x"F2B4",
		x"F2B5", x"F1D7", x"F001", x"EDA5", x"EBEF", x"EC1E", x"EF35", x"F53A",
		x"FD2D", x"05C6", x"0D48", x"124B", x"1403", x"1286", x"0E95", x"090B",
		x"02C8", x"FC63", x"F6A1", x"F1E8", x"EE95", x"EC87", x"EB4F", x"EAD0",
		x"EAB8", x"EAF4", x"EBA2", x"ED1A", x"F022", x"F501", x"FB86", x"02FD",
		x"0A2F", x"0FFF", x"137C", x"148D", x"1389", x"1150", x"0EBA", x"0C10",
		x"0A44", x"09E1", x"0B38", x"0DD4", x"10CF", x"12B4", x"1267", x"0F29",
		x"0952", x"027E", x"FCA7", x"F9BA", x"FAA2", x"FF2F", x"05D6", x"0C80",
		x"113A", x"12E0", x"11A8", x"0ECE", x"0BB1", x"09A1", x"0977", x"0AED",
		x"0D6C", x"101C", x"126B", x"13D3", x"13EE", x"1237", x"0E6A", x"0897",
		x"013D", x"F982", x"F2A7", x"EDDD", x"EB88", x"EB36", x"EC03", x"ED27",
		x"EE62", x"EF6E", x"F08E", x"F1A8", x"F30B", x"F529", x"F7FA", x"FBA1",
		x"FF90", x"0360", x"0678", x"0846", x"08E1", x"082B", x"0691", x"03F9",
		x"00C2", x"FD1E", x"F9A9", x"F712", x"F5DB", x"F697", x"F99F", x"FEC5",
		x"0527", x"0BA1", x"10D2", x"1341", x"1267", x"0E2B", x"0787", x"FFEE",
		x"F88F", x"F253", x"EDF2", x"EBBE", x"EBFE", x"EF2F", x"F4FF", x"FCD3",
		x"0555", x"0CD7", x"120C", x"1440", x"13EE", x"1211", x"0FE9", x"0E80",
		x"0E40", x"0F10", x"1063", x"11CC", x"131E", x"1433", x"14D5", x"14BD",
		x"13B5", x"11A4", x"0EBD", x"0B6A", x"08B9", x"079B", x"0888", x"0B5C",
		x"0EFF", x"11F7", x"12E3", x"10E4", x"0BEB", x"0561", x"FF6A", x"FC1C",
		x"FC7D", x"0062", x"0665", x"0CB2", x"1130", x"129A", x"10BC", x"0C33",
		x"0678", x"00BE", x"FBCE", x"F804", x"F548", x"F3CF", x"F389", x"F498",
		x"F723", x"FBA1", x"01D8", x"08D2", x"0EC7", x"1270", x"136A", x"11FB",
		x"0F9F", x"0DBD", x"0D82", x"0EDF", x"1101", x"1305", x"146C", x"153A",
		x"158C", x"156A", x"1520", x"14A5", x"137F", x"1181", x"0F4F", x"0DC8",
		x"0DE0", x"0F75", x"1188", x"12E8", x"1252", x"0F2C", x"0987", x"0245",
		x"FB58", x"F631", x"F38B", x"F320", x"F441", x"F68B", x"F9BA", x"FDD6",
		x"0251", x"06A7", x"0A26", x"0CB8", x"0E97", x"0FEA", x"112E", x"1261",
		x"1358", x"142C", x"148D", x"14B5", x"1476", x"13C0", x"1285", x"1108",
		x"0F67", x"0E5E", x"0E4B", x"0F28", x"10AA", x"1244", x"136E", x"146F",
		x"1508", x"151F", x"14E8", x"14B3", x"14C2", x"14E3", x"1528", x"14F8",
		x"143A", x"12AD", x"0FF9", x"0B64", x"04DC", x"FCCC", x"F4F4", x"EF0E",
		x"EC4A", x"EC0C", x"ED34", x"EE22", x"EE09", x"ED22", x"ECB1", x"EE4A",
		x"F2C9", x"F9F1", x"0226", x"0989", x"0F07", x"1268", x"1429", x"14EB",
		x"151F", x"1525", x"1518", x"14FF", x"14A6", x"1400", x"1321", x"120E",
		x"10F3", x"0F67", x"0D02", x"099F", x"0502", x"FF36", x"F8BA", x"F268",
		x"EDF5", x"EC8A", x"EE44", x"F1E5", x"F5BF", x"F83B", x"F863", x"F67E",
		x"F363", x"F035", x"ED98", x"EBDA", x"EB15", x"EBD4", x"EF2C", x"F568",
		x"FDA8", x"0627", x"0D62", x"1245", x"1503", x"15DC", x"1508", x"1295",
		x"0DF4", x"073B", x"FF18", x"F6EF", x"F052", x"EC6F", x"EBF5", x"EEAC",
		x"F437", x"FB8F", x"03D3", x"0B8C", x"1179", x"14CD", x"15A3", x"1538",
		x"14B5", x"1499", x"1493", x"1441", x"132C", x"1166", x"0F1A", x"0CA1",
		x"0A40", x"0821", x"0660", x"048B", x"0255", x"FFD0", x"FCEF", x"F9CA",
		x"F684", x"F362", x"F0B3", x"EE9D", x"ED27", x"EC54", x"EBF3", x"EC19",
		x"EC77", x"ED22", x"EE14", x"EF6C", x"F150", x"F39E", x"F651", x"F98A",
		x"FD7E", x"0204", x"0669", x"0A22", x"0CE4", x"0E9F", x"0F31", x"0E28",
		x"0ADE", x"052B", x"FDBD", x"F60B", x"EFFC", x"ECB8", x"EC1D", x"ECEB",
		x"ED8D", x"ED48", x"EC97", x"ED1D", x"F037", x"F647", x"FE92", x"0700",
		x"0DD6", x"1231", x"1426", x"14D4", x"14D4", x"14C4", x"14BA", x"14A4",
		x"1407", x"11D7", x"0DB1", x"0748", x"FFA3", x"F7FE", x"F1A9", x"ED39",
		x"EB2A", x"EB4D", x"ED33", x"F01D", x"F365", x"F631", x"F89B", x"FA67",
		x"FB33", x"FAED", x"F98A", x"F713", x"F404", x"F10A", x"EE81", x"ECD0",
		x"EC06", x"EC60", x"EE6E", x"F2F0", x"F9CE", x"01E4", x"09A9", x"0FB0",
		x"135E", x"151C", x"15AE", x"157A", x"1455", x"118E", x"0C73", x"04FF",
		x"FC68", x"F458", x"EEDD", x"ECCB", x"EE51", x"F29D", x"F8D0", x"FFC8",
		x"06CB", x"0C98", x"10EB", x"1394", x"14C4", x"14DC", x"1427", x"1317",
		x"1216", x"116C", x"113E", x"118B", x"1241", x"1349", x"1471", x"151E",
		x"151F", x"14C8", x"144C", x"1457", x"14B8", x"1525", x"1527", x"148D",
		x"136C", x"1231", x"1194", x"11AA", x"129D", x"13AB", x"13DF", x"1233",
		x"0E01", x"074F", x"FEFD", x"F6C6", x"F050", x"ED0A", x"ED75", x"F140",
		x"F770", x"FE80", x"052F", x"0A8D", x"0DF3", x"0F67", x"0F09", x"0D69",
		x"0AD8", x"07E5", x"04A2", x"01B7", x"FF86", x"FE7E", x"FEC1", x"0043",
		x"02A7", x"059D", x"08B4", x"0BB6", x"0E86", x"10DB", x"12E9", x"1422",
		x"14A0", x"1483", x"1413", x"13E4", x"1432", x"14C7", x"1500", x"13DE",
		x"108E", x"0AE4", x"0346", x"FB0F", x"F3E9", x"EF12", x"ECD2", x"ECAE",
		x"EE0C", x"F051", x"F39D", x"F782", x"FB06", x"FD3C", x"FDA7", x"FC51",
		x"F97A", x"F604", x"F278", x"EF97", x"EDC0", x"ED2E", x"EDED", x"F058",
		x"F4F0", x"FB81", x"0313", x"0A6F", x"102E", x"137F", x"144D", x"12AB",
		x"0F8A", x"0BFA", x"08DC", x"068A", x"04FC", x"0411", x"03A1", x"03D6",
		x"048A", x"05A6", x"0753", x"0974", x"0BC1", x"0E18", x"103D", x"11FF",
		x"1363", x"143C", x"1480", x"1404", x"1352", x"12BC", x"125C", x"1247",
		x"1291", x"134C", x"1445", x"1508", x"150A", x"1481", x"13C3", x"13B7",
		x"1432", x"14A1", x"1400", x"1169", x"0C36", x"04C2", x"FC83", x"F510",
		x"EFA3", x"EC80", x"EB42", x"EB6E", x"EC50", x"ED58", x"EDEC", x"EDE1",
		x"ED1E", x"EC3A", x"EBB9", x"ECBB", x"F012", x"F5F1", x"FD94", x"0565",
		x"0C21", x"10EC", x"13B1", x"14FA", x"1560", x"1549", x"14FF", x"14A1",
		x"1439", x"136C", x"11DB", x"0F5D", x"0C17", x"0829", x"0492", x"01E0",
		x"00D7", x"01BF", x"04C7", x"0969", x"0E72", x"1230", x"1327", x"10E9",
		x"0C37", x"0640", x"0069", x"FBAC", x"F86E", x"F693", x"F57B", x"F428",
		x"F250", x"F021", x"EDAD", x"EC12", x"EBE9", x"ED8F", x"F170", x"F77F",
		x"FF50", x"076E", x"0E6B", x"12B6", x"138E", x"10E2", x"0B41", x"03E4",
		x"FC61", x"F5FC", x"F161", x"EEFB", x"EEA8", x"EFE0", x"F24C", x"F583",
		x"F901", x"FC28", x"FE10", x"FDF3", x"FB9E", x"F783", x"F29C", x"EE7A",
		x"ECF8", x"EED8", x"F409", x"FB7A", x"0384", x"0AF0", x"1075", x"13BF",
		x"14AA", x"1314", x"0EE6", x"0835", x"0014", x"F7EE", x"F141", x"ED6B",
		x"ECEE", x"EF75", x"F3AC", x"F801", x"FB3F", x"FCCB", x"FC76", x"FA89",
		x"F7C8", x"F4DF", x"F21D", x"EFE4", x"EE66", x"ED9D", x"EDA3", x"EE47",
		x"EF50", x"F0D5", x"F337", x"F69D", x"FB68", x"0190", x"085E", x"0E93",
		x"12BF", x"13B5", x"1162", x"0CF7", x"087C", x"061B", x"069B", x"09F0",
		x"0E77", x"1214", x"130A", x"106C", x"0B00", x"03FC", x"FD3A", x"F795",
		x"F381", x"F104", x"EF90", x"EE9F", x"EDE9", x"EDA8", x"EDC1", x"EEB0",
		x"F07C", x"F2FE", x"F609", x"F91D", x"FB96", x"FC85", x"FB9F", x"F898",
		x"F42A", x"EFB5", x"ED40", x"EE11", x"F259", x"F86B", x"FDDC", x"00DD",
		x"00DD", x"FE6F", x"FAB2", x"F6AB", x"F302", x"F04E", x"EF27", x"F042",
		x"F459", x"FB04", x"0342", x"0B20", x"10E8", x"13BF", x"1405", x"12E7",
		x"11E2", x"11DA", x"12D1", x"13F4", x"14B9", x"14C4", x"1469", x"13E2",
		x"13BC", x"1402", x"147D", x"14C7", x"149F", x"13FD", x"130D", x"124C",
		x"11C1", x"11CA", x"1272", x"1376", x"14A5", x"154B", x"1570", x"14FA",
		x"140B", x"12DA", x"114A", x"0F9E", x"0DBF", x"0BED", x"09C5", x"0765",
		x"04AF", x"01CC", x"FEFB", x"FC71", x"FA1D", x"F7E6", x"F5BD", x"F395",
		x"F17F", x"EF71", x"EDA8", x"EC56", x"EB72", x"EB0F", x"EAD9", x"EAE4",
		x"EB12", x"EB5C", x"EB99", x"EBBE", x"EB9E", x"EB7E", x"EB8F", x"EC09",
		x"ED5C", x"EFEA", x"F3CD", x"F934", x"FF9E", x"06A7", x"0D09", x"11A2",
		x"139F", x"129E", x"0EBB", x"088B", x"011C", x"F984", x"F310", x"EE8B",
		x"EC58", x"ECB2", x"EFC8", x"F566", x"FCDE", x"04F0", x"0BF1", x"1109",
		x"138F", x"13BA", x"120A", x"0F7F", x"0CDC", x"0A60", x"0873", x"071F",
		x"05B3", x"0374", x"FFA8", x"FA51", x"F46A", x"EF94", x"ED73", x"EF04",
		x"F3B2", x"F9A0", x"FE93", x"0088", x"FE9C", x"F992", x"F33F", x"EE2A",
		x"EC8E", x"EE5D", x"F20E", x"F56E", x"F6AE", x"F546", x"F228", x"EEA3",
		x"ECC6", x"EE3E", x"F38E", x"FBE5", x"0543", x"0D71", x"126D", x"138D",
		x"1115", x"0C3E", x"06CF", x"0253", x"0030", x"0124", x"04E4", x"0A30",
		x"0F52", x"1293", x"12B3", x"0F77", x"09C1", x"0328", x"FD6D", x"F92A",
		x"F64E", x"F498", x"F393", x"F303", x"F2BA", x"F2B0", x"F2CB", x"F359",
		x"F43B", x"F599", x"F7DF", x"FB53", x"FFF0", x"0579", x"0B35", x"1041",
		x"1385", x"1416", x"118A", x"0C4C", x"05B8", x"FF4F", x"FA1B", x"F63B",
		x"F37D", x"F1A2", x"F05B", x"EF59", x"EE2F", x"ECA3", x"EB77", x"EBEA",
		x"EEF7", x"F4BF", x"FC71", x"04AC", x"0C0A", x"115D", x"1459", x"1501",
		x"140B", x"11F6", x"0F14", x"0BC6", x"08BD", x"06C1", x"06E2", x"094E",
		x"0D3F", x"10F3", x"1272", x"109C", x"0BCC", x"05B2", x"008B", x"FE2F",
		x"FF93", x"03FF", x"09FF", x"0F8E", x"12DC", x"12BA", x"0EFC", x"0830",
		x"FF9A", x"F71C", x"F06D", x"ECA4", x"EBE3", x"ED7E", x"F0C4", x"F529",
		x"F9E4", x"FE4C", x"01D1", x"0493", x"06E5", x"08F8", x"0AB4", x"0C5E",
		x"0E01", x"0FB5", x"114F", x"127A", x"134E", x"1404", x"14A3", x"150B",
		x"14F0", x"140D", x"124F", x"0FE4", x"0D40", x"0ACB", x"0917", x"0891",
		x"0995", x"0BE4", x"0F0E", x"1217", x"1403", x"13A2", x"1041", x"09FD",
		x"01A5", x"F8F9", x"F1E5", x"EDF0", x"EDF7", x"F185", x"F73F", x"FD5E",
		x"01E4", x"0376", x"014E", x"FC01", x"F545", x"EFC3", x"ED42", x"EE05",
		x"F0BC", x"F347", x"F424", x"F2CB", x"F002", x"EDA4", x"EDA8", x"F12B",
		x"F7BD", x"FF78", x"06E0", x"0CB0", x"10BC", x"132E", x"1472", x"14CB",
		x"14CE", x"14A3", x"1406", x"1236", x"0E81", x"08A2", x"011A", x"F913",
		x"F206", x"ED27", x"EAB1", x"EA36", x"EA8C", x"EAE0", x"EB00", x"EBA1",
		x"ECF9", x"EEFC", x"F19D", x"F476", x"F6FE", x"F8B1", x"F9BB", x"FA90",
		x"FC0A", x"FEC9", x"02E6", x"07DB", x"0CD8", x"10CB", x"12BC", x"11EF",
		x"0E6C", x"08D8", x"02A1", x"FD3E", x"F9AB", x"F84D", x"F8B7", x"FAC2",
		x"FE2B", x"0267", x"06BE", x"0AA0", x"0D86", x"0F88", x"10D7", x"11B3",
		x"1262", x"131A", x"13E1", x"1491", x"147B", x"1277", x"0D62", x"05A7",
		x"FCB9", x"F4D2", x"EF31", x"EC00", x"EAAF", x"EAD3", x"ECD5", x"F0D4",
		x"F6E2", x"FE7D", x"067A", x"0D78", x"124C", x"149A", x"154F", x"1552",
		x"151E", x"14D3", x"13D6", x"11A8", x"0DE6", x"0867", x"016D", x"F9D9",
		x"F2EF", x"EE1E", x"EC58", x"ED48", x"EF91", x"F186", x"F1F6", x"F075",
		x"EE2D", x"ED3F", x"EF38", x"F49B", x"FBF4", x"02F0", x"07CE", x"09B4",
		x"08CD", x"05D7", x"01CA", x"FD3A", x"F8E3", x"F5AC", x"F42D", x"F4D9",
		x"F778", x"FB2E", x"FF75", x"037D", x"06AE", x"0826", x"07B4", x"0504",
		x"004C", x"FA1F", x"F3BD", x"EED1", x"EC99", x"ED5E", x"F078", x"F4FF",
		x"F9F5", x"FEB0", x"02B0", x"05E7", x"0828", x"099A", x"0A29", x"09D3",
		x"08EC", x"0732", x"04EF", x"01F6", x"FECB", x"FB95", x"F8FE", x"F786",
		x"F750", x"F893", x"FAFE", x"FE67", x"0230", x"05BB", x"088B", x"0A29",
		x"0A87", x"093E", x"0677", x"02A8", x"FE67", x"FA92", x"F7E3", x"F6FC",
		x"F812", x"FB74", x"0107", x"0790", x"0DBF", x"11EB", x"133A", x"11C0",
		x"0E3D", x"0982", x"04A1", x"0073", x"FD27", x"FAA8", x"F8F9", x"F7E6",
		x"F782", x"F7B1", x"F83F", x"F96E", x"FB41", x"FDDA", x"00F2", x"044E",
		x"0780", x"0A72", x"0D1B", x"0F38", x"10D6", x"11F7", x"12E7", x"1389",
		x"142C", x"148D", x"1483", x"13DD", x"128E", x"1074", x"0E52", x"0C76",
		x"0B7C", x"0BDD", x"0D8E", x"101B", x"1294", x"13AE", x"1254", x"0E42",
		x"07F8", x"0094", x"F959", x"F35E", x"EF22", x"EC85", x"EB42", x"EAE8",
		x"EAD8", x"EADF", x"EB2F", x"EC0A", x"EE0A", x"F1AA", x"F758", x"FEC5",
		x"06EE", x"0DFD", x"1283", x"1399", x"1137", x"0BE9", x"04C0", x"FD48",
		x"F68C", x"F13D", x"EDB9", x"EBEE", x"EBDA", x"ED58", x"EF92", x"F212",
		x"F461", x"F5D5", x"F5F1", x"F48A", x"F1FD", x"EF05", x"ECDD", x"EC99",
		x"EEFC", x"F42E", x"FB5D", x"02BE", x"08F8", x"0D54", x"0FD5", x"1126",
		x"11CB", x"1275", x"1354", x"146E", x"14E8", x"13BC", x"0FE1", x"0932",
		x"00D0", x"F88F", x"F1E2", x"ED85", x"EB54", x"EB7E", x"EE01", x"F2B6",
		x"F96F", x"0166", x"0945", x"0FAC", x"138B", x"1545", x"1578", x"154B",
		x"1537", x"14EF", x"1406", x"1225", x"0EFF", x"0ABA", x"0570", x"FF65",
		x"F91E", x"F325", x"EE98", x"EC3E", x"ECE4", x"F0B3", x"F739", x"FF70",
		x"07D5", x"0EC1", x"1312", x"147F", x"139B", x"110F", x"0D89", x"097C",
		x"050B", x"00FB", x"FD48", x"FA7A", x"F8B7", x"F81E", x"F8AE", x"FA7A",
		x"FD4D", x"00DE", x"04C5", x"0819", x"0A60", x"0B33", x"0A8B", x"084B",
		x"0469", x"FF12", x"F8DF", x"F2BC", x"EE4E", x"ECCF", x"EF1A", x"F513",
		x"FD91", x"0675", x"0E06", x"12DE", x"1457", x"1366", x"11B0", x"10DB",
		x"1177", x"12D6", x"1371", x"11A1", x"0CE3", x"05A9", x"FDC5", x"F735",
		x"F36C", x"F27F", x"F401", x"F70C", x"FB64", x"0035", x"0494", x"0768",
		x"083C", x"06D4", x"0399", x"FF66", x"FABC", x"F6AB", x"F3D5", x"F2D3",
		x"F42E", x"F822", x"FE71", x"05FF", x"0D17", x"11F4", x"13DC", x"1363",
		x"116E", x"0F65", x"0E4D", x"0E72", x"0FBB", x"118F", x"135F", x"146E",
		x"14D0", x"1448", x"1327", x"11AD", x"1016", x"0E4F", x"0C6F", x"0ACE",
		x"098F", x"091A", x"09B5", x"0B1F", x"0D2A", x"0F67", x"1165", x"12FA",
		x"141C", x"14B7", x"14CB", x"144E", x"1353", x"11F5", x"0FEE", x"0DAF",
		x"0B5F", x"0996", x"087E", x"0858", x"0907", x"0A42", x"0BFC", x"0E14",
		x"108A", x"12D5", x"145F", x"141C", x"11A5", x"0C92", x"0581", x"FD8B",
		x"F61A", x"F07B", x"ED1C", x"EBC6", x"EB9F", x"EC2C", x"ED36", x"EEB6",
		x"F101", x"F402", x"F74B", x"FA70", x"FD4C", x"FFD8", x"0251", x"04DF",
		x"079A", x"0A48", x"0CBB", x"0E94", x"0FDF", x"10DC", x"11BC", x"129E",
		x"1378", x"143B", x"149E", x"1425", x"1219", x"0DD4", x"0762", x"FFA2",
		x"F7FD", x"F1AB", x"ED83", x"EB98", x"EB2C", x"EB4C", x"EB63", x"EB29",
		x"EADB", x"EAFC", x"EC01", x"EE49", x"F261", x"F891", x"003E", x"083C",
		x"0ED3", x"12BE", x"1423", x"13CF", x"1302", x"12B4", x"134A", x"1406",
		x"13B9", x"10F8", x"0B17", x"02CF", x"F9C8", x"F22F", x"EDC3", x"ED38",
		x"F03A", x"F586", x"FBDF", x"01EA", x"070E", x"0B03", x"0D66", x"0EA8",
		x"0EA1", x"0D76", x"0B19", x"073F", x"023D", x"FC66", x"F685", x"F15C",
		x"EDA4", x"EC02", x"ECFD", x"F080", x"F603", x"FC83", x"0308", x"08FF",
		x"0DCF", x"114A", x"1353", x"1449", x"1464", x"13CB", x"126B", x"0FDA",
		x"0BDD", x"0641", x"FF86", x"F857", x"F201", x"EDBB", x"EC2D", x"ED2A",
		x"EFD4", x"F341", x"F6BF", x"F983", x"FB10", x"FB11", x"F98E", x"F70B",
		x"F3E0", x"F073", x"ED9B", x"EC65", x"EDC6", x"F229", x"F930", x"01BE",
		x"09E6", x"1025", x"1341", x"1305", x"1043", x"0BBA", x"066A", x"00FB",
		x"FC26", x"F823", x"F522", x"F333", x"F1C4", x"F069", x"EED0", x"ECFB",
		x"EBBB", x"EB9B", x"ED84", x"F1D9", x"F852", x"0041", x"080B", x"0E92",
		x"12C4", x"14D5", x"1542", x"1517", x"1513", x"1504", x"14C8", x"13E5",
		x"11BF", x"0D70", x"0688", x"FDCD", x"F532", x"EEEB", x"EBF9", x"EB83",
		x"EC21", x"EC7A", x"EC7C", x"ECCB", x"EEE2", x"F38D", x"FAA2", x"029B",
		x"097B", x"0D58", x"0D8A", x"0A51", x"047D", x"FD30", x"F5CA", x"EFFC",
		x"ED3F", x"EE96", x"F373", x"FA6A", x"01D7", x"08A9", x"0E52", x"126F",
		x"1437", x"131F", x"0F0E", x"08BD", x"00F4", x"F91A", x"F248", x"ED7C",
		x"EB73", x"EBF3", x"EE42", x"F14B", x"F4B5", x"F7BE", x"FA7F", x"FCE6",
		x"FEB7", x"FFE5", x"007F", x"0085", x"FFE1", x"FEB8", x"FCDF", x"FA8B",
		x"F7D7", x"F4ED", x"F1A3", x"EE89", x"EC47", x"EBBB", x"EDB7", x"F24C",
		x"F8D3", x"00A1", x"0879", x"0F10", x"1334", x"145A", x"129F", x"0E7C",
		x"0870", x"0131", x"F9D3", x"F334", x"EE7F", x"ECD1", x"EE91", x"F39C",
		x"FA9F", x"01FC", x"0862", x"0CF5", x"0F7A", x"1004", x"0EDB", x"0C29",
		x"0872", x"0442", x"00C8", x"FF07", x"FFD6", x"035F", x"08D6", x"0E84",
		x"11F5", x"11BF", x"0E3E", x"096A", x"060B", x"05E7", x"0925", x"0E0A",
		x"1201", x"12AD", x"0FA5", x"0A63", x"0554", x"02E3", x"0415", x"0863",
		x"0DDF", x"1232", x"1358", x"10C8", x"0B58", x"0482", x"FDF1", x"F88A",
		x"F4E4", x"F2BA", x"F1B2", x"F112", x"F07A", x"EFF9", x"EFBA", x"F01C",
		x"F131", x"F2DB", x"F4E6", x"F75C", x"FA56", x"FDDE", x"01AC", x"0557",
		x"08A0", x"0B7F", x"0DED", x"0FB0", x"10BA", x"114C", x"1178", x"1194",
		x"117C", x"110E", x"1023", x"0E71", x"0BC7", x"07D1", x"029F", x"FC50",
		x"F5C0", x"F01B", x"ECD3", x"ECD7", x"EFF5", x"F4BC", x"F979", x"FC97",
		x"FD7B", x"FC21", x"F93E", x"F5EE", x"F2CD", x"F06E", x"EEDD", x"EED7",
		x"F0AC", x"F500", x"FB90", x"0355", x"0AD4", x"1065", x"135C", x"13B4",
		x"11FE", x"0F82", x"0D54", x"0BF8", x"0B1C", x"09DA", x"0790", x"03BF",
		x"FE82", x"F868", x"F2A4", x"EE7C", x"ED10", x"EEB2", x"F2B8", x"F79F",
		x"FC23", x"FEAA", x"FF4A", x"FE02", x"FB50", x"F7C8", x"F41E", x"F0E5",
		x"EE73", x"ECD2", x"EBC9", x"EB57", x"EB33", x"EB1C", x"EB29", x"EB50",
		x"EC3B", x"EE7D", x"F2B0", x"F8CA", x"0030", x"07E2", x"0E5A", x"12A7",
		x"1413", x"128F", x"0E21", x"0740", x"FF33", x"F75C", x"F13D", x"ED67",
		x"EBE6", x"EC43", x"EDD9", x"F008", x"F21A", x"F391", x"F4B3", x"F612",
		x"F85F", x"FBEF", x"010E", x"073E", x"0D58", x"1198", x"12CD", x"1086",
		x"0BEF", x"0763", x"0536", x"068E", x"0A9B", x"0F37", x"11D2", x"10F4",
		x"0CCA", x"074E", x"034F", x"02D8", x"0657", x"0BEB", x"10D2", x"127F",
		x"1015", x"0B4A", x"06D5", x"0540", x"0739", x"0BCD", x"106F", x"126B",
		x"108B", x"0B9D", x"0627", x"02E1", x"0348", x"0702", x"0C42", x"10C4",
		x"128B", x"1103", x"0CB3", x"06DE", x"00B9", x"FB2B", x"F6C3", x"F3C4",
		x"F1E2", x"F0F1", x"F090", x"F066", x"F07F", x"F0EF", x"F1BB", x"F32E",
		x"F549", x"F7D3", x"FAD2", x"FDF5", x"0144", x"046E", x"0744", x"09E1",
		x"0C24", x"0E1D", x"0FE8", x"113C", x"1247", x"134F", x"1442", x"14EB",
		x"154D", x"1546", x"1509", x"1448", x"127F", x"0F15", x"09A9", x"0260",
		x"FA4A", x"F340", x"EE59", x"EC43", x"EC15", x"ECCC", x"ED48", x"ED40",
		x"ECA7", x"EBB1", x"EAFA", x"EAC4", x"EAED", x"EB2E", x"EB49", x"EBA0",
		x"ED0C", x"F084", x"F692", x"FEA4", x"071E", x"0E6D", x"1334", x"14B2",
		x"12F9", x"0E98", x"086C", x"015B", x"FA3F", x"F3C4", x"EED3", x"EC95",
		x"EDC6", x"F24E", x"F916", x"00AF", x"07BA", x"0D33", x"10F3", x"12D7",
		x"136B", x"12FF", x"11D6", x"0FC4", x"0CD1", x"091B", x"054A", x"01FB",
		x"FF5E", x"FD89", x"FC4D", x"FB0E", x"F980", x"F724", x"F3E3", x"F06D",
		x"EDBC", x"ED46", x"EFC9", x"F51F", x"FC34", x"036A", x"0926", x"0C70",
		x"0C8F", x"098A", x"03E1", x"FC97", x"F52D", x"EF5F", x"EC68", x"ECBF",
		x"EFC3", x"F45A", x"F973", x"FE17", x"01BB", x"0421", x"0502", x"044B",
		x"01C6", x"FD62", x"F77E", x"F1B4", x"EDC8", x"ECEB", x"EF36", x"F31C",
		x"F680", x"F74C", x"F50E", x"F0F5", x"EDA0", x"ED74", x"F12C", x"F773",
		x"FDFB", x"029C", x"0406", x"027E", x"FEB1", x"FA26", x"F5CA", x"F29D",
		x"F104", x"F17B", x"F4B4", x"FAA1", x"0284", x"0A72", x"108C", x"13BB",
		x"143E", x"1309", x"1140", x"101F", x"1044", x"118C", x"1359", x"14BE",
		x"1571", x"1578", x"14C8", x"1351", x"1127", x"0EC8", x"0C54", x"0A2D",
		x"0860", x"073E", x"06F6", x"079F", x"0918", x"0AF8", x"0D32", x"0F6C",
		x"1175", x"12FD", x"1409", x"1464", x"1419", x"132E", x"11BC", x"0FB3",
		x"0D26", x"0A37", x"071C", x"0453", x"01F6", x"0024", x"FEAB", x"FD4F",
		x"FB64", x"F893", x"F4EF", x"F103", x"EDC5", x"EC49", x"ED80", x"F175",
		x"F7D2", x"FF20", x"0600", x"0AFD", x"0DC7", x"0E88", x"0DB3", x"0B7D",
		x"083C", x"0441", x"0038", x"FC63", x"F91E", x"F67A", x"F48F", x"F333",
		x"F1DB", x"F073", x"EE93", x"ECCD", x"EBAD", x"EB86", x"ED1B", x"F097",
		x"F63F", x"FD59", x"0542", x"0C6E", x"118F", x"13B1", x"121E", x"0D11",
		x"05E4", x"FE11", x"F707", x"F1B0", x"EE59", x"EC74", x"EB94", x"EB60",
		x"EB8F", x"EC56", x"EE10", x"F0B9", x"F4B5", x"FA3E", x"012D", x"08B6",
		x"0F2A", x"1305", x"1367", x"10F5", x"0DA0", x"0B7A", x"0B93", x"0DE7",
		x"10F0", x"127B", x"10C4", x"0B86", x"04AA", x"FED5", x"FC79", x"FE72",
		x"03FF", x"0ACE", x"1038", x"128B", x"1141", x"0DD8", x"0A29", x"0811",
		x"083E", x"0A7D", x"0DEA", x"1118", x"1346", x"147E", x"14BD", x"13B7",
		x"10EE", x"0BE7", x"04F7", x"FD04", x"F594", x"EFC0", x"EC65", x"EB7A",
		x"EC6A", x"EE76", x"F0EC", x"F347", x"F506", x"F61B", x"F691", x"F696",
		x"F62A", x"F544", x"F3D3", x"F220", x"F04E", x"EE96", x"ED02", x"EBB3",
		x"EAD5", x"EAAD", x"EB3F", x"EC6D", x"EDDD", x"EF0C", x"EFF3", x"F0AE",
		x"F118", x"F121", x"F0CE", x"F026", x"EF19", x"EDCD", x"EC40", x"EB2E",
		x"EB90", x"EDF9", x"F269", x"F89E", x"FFFF", x"076D", x"0DD3", x"1234",
		x"1466", x"148E", x"132D", x"10D5", x"0DF3", x"0B1B", x"091F", x"087E",
		x"094C", x"0B9C", x"0ECE", x"11EE", x"139C", x"12B7", x"0ED2", x"08A1",
		x"019D", x"FB08", x"F5F8", x"F296", x"F083", x"EF52", x"EE9A", x"EDC2",
		x"ECAD", x"EBAB", x"EBAE", x"EE54", x"F408", x"FBE0", x"0434", x"0B91",
		x"1106", x"1422", x"14DA", x"1318", x"0F30", x"093A", x"01A7", x"F957",
		x"F209", x"ED10", x"EB02", x"EB20", x"EC64", x"EDC8", x"EEDA", x"EFD9",
		x"F136", x"F354", x"F69B", x"FAF8", x"009E", x"06FA", x"0D16", x"11BF",
		x"13CB", x"1289", x"0DEF", x"0722", x"FF3B", x"F791", x"F132", x"ECEA",
		x"EB63", x"EC64", x"EF86", x"F3E9", x"F905", x"FE58", x"0378", x"07C0",
		x"0ACA", x"0C59", x"0C6B", x"0AC7", x"0701", x"00EC", x"F949", x"F239",
		x"ED9C", x"EC32", x"ED70", x"EF78", x"F0AB", x"F00E", x"EE38", x"EC75",
		x"EC92", x"EFCF", x"F663", x"FF5F", x"089B", x"0FAA", x"12F3", x"11EF",
		x"0D95", x"0762", x"00D4", x"FB76", x"F86F", x"F92A", x"FD55", x"03EB",
		x"0ACE", x"100A", x"12B1", x"1279", x"1067", x"0DA5", x"0BD1", x"0B6E",
		x"0C85", x"0EC3", x"113B", x"135B", x"14A9", x"14FF", x"1486", x"1344",
		x"117B", x"0F54", x"0D50", x"0BF1", x"0B6F", x"0C25", x"0E06", x"10AF",
		x"12DF", x"1341", x"10DE", x"0B91", x"044C", x"FCC7", x"F671", x"F1FF",
		x"EF39", x"EDB6", x"ECB2", x"EBF5", x"EB7B", x"EB1E", x"EAF0", x"EB0B",
		x"EBC1", x"ED3A", x"EFA5", x"F253", x"F467", x"F50E", x"F420", x"F1DA",
		x"EF29", x"ED42", x"EDA6", x"F10C", x"F743", x"FE71", x"049F", x"0861",
		x"096F", x"080C", x"04D7", x"0098", x"FC6B", x"F93F", x"F7BB", x"F802",
		x"FA4B", x"FE9C", x"0493", x"0B27", x"10A8", x"13A5", x"12E8", x"0E78",
		x"0731", x"FE9F", x"F662", x"F015", x"ECA9", x"EBFD", x"ED62", x"EFCD",
		x"F206", x"F32D", x"F2CD", x"F147", x"EF2D", x"ED36", x"EBD6", x"EB34",
		x"EB03", x"EAFC", x"EAFC", x"EB46", x"EC11", x"ED64", x"EF46", x"F174",
		x"F3C2", x"F5E4", x"F7C5", x"F947", x"FAD8", x"FCBB", x"FF37", x"02BF",
		x"071F", x"0BEF", x"105A", x"1323", x"1378", x"10C9", x"0B59", x"0467",
		x"FDE0", x"F964", x"F78E", x"F816", x"FA2F", x"FD76", x"017D", x"058E",
		x"08EC", x"0AD7", x"0AEE", x"0943", x"063B", x"027F", x"FEA0", x"FB4C",
		x"F91C", x"F8A5", x"FA23", x"FDC1", x"0317", x"0941", x"0EFF", x"12C1",
		x"1383", x"10A0", x"0A63", x"0213", x"F961", x"F225", x"ED80", x"EBF4",
		x"ECEA", x"EF73", x"F24C", x"F47A", x"F55D", x"F4E2", x"F350", x"F119",
		x"EED4", x"ED0C", x"EBE6", x"EB43", x"EB4A", x"EBE3", x"ED0E", x"EEA4",
		x"F050", x"F191", x"F231", x"F244", x"F177", x"EFE0", x"EDFA", x"EC4E",
		x"EB69", x"EB28", x"EB0F", x"EAD1", x"EB3A", x"ED1A", x"F184", x"F81A",
		x"003B", x"087D", x"0F55", x"13B3", x"159F", x"159A", x"1462", x"1288",
		x"101E", x"0D48", x"0A9F", x"093B", x"09DE", x"0C73", x"0FF9", x"1274",
		x"1251", x"0F0F", x"094B", x"02BE", x"FD30", x"F9C0", x"F890", x"F939",
		x"FB6A", x"FEB5", x"029F", x"06B1", x"0A8A", x"0DCE", x"1054", x"1224",
		x"136E", x"143B", x"14B7", x"14E7", x"150F", x"152C", x"1546", x"1549",
		x"1514", x"1483", x"137C", x"1215", x"1050", x"0E38", x"0BE1", x"095A",
		x"06E4", x"047D", x"020B", x"FF82", x"FCEA", x"FA6B", x"F826", x"F62D",
		x"F495", x"F32C", x"F1BA", x"F023", x"EE5E", x"ECB5", x"EB8E", x"EBED",
		x"EE61", x"F37B", x"FAA2", x"029A", x"09F4", x"0F86", x"1309", x"14A1",
		x"1519", x"14F3", x"143E", x"12EC", x"10B0", x"0D76", x"0933", x"03EF",
		x"FE0C", x"F7D8", x"F249", x"EE04", x"EC10", x"ED1F", x"F145", x"F7DE",
		x"FF7F", x"0704", x"0D4C", x"11C8", x"13F8", x"1368", x"1019", x"0A72",
		x"0313", x"FB25", x"F3F0", x"EECC", x"EC82", x"ED03", x"EF94", x"F310",
		x"F627", x"F824", x"F8B6", x"F7E8", x"F60D", x"F362", x"F063", x"EDC0",
		x"EBF9", x"EBCA", x"ED6A", x"F101", x"F667", x"FD20", x"0475", x"0B37",
		x"1080", x"12C5", x"113E", x"0BE9", x"03F5", x"FB68", x"F456", x"EFA1",
		x"ED64", x"ECFD", x"EEA2", x"F24E", x"F815", x"FF75", x"075F", x"0E31",
		x"1282", x"13D6", x"1279", x"0F9E", x"0C55", x"0965", x"076A", x"0684",
		x"06E2", x"0871", x"0AF1", x"0E43", x"119B", x"13D5", x"13E4", x"111E",
		x"0B54", x"035D", x"FA95", x"F2C0", x"EDB1", x"EC41", x"EE29", x"F240",
		x"F71B", x"FBC1", x"FF77", x"0222", x"03AF", x"0423", x"0344", x"00D1",
		x"FCBB", x"F7A8", x"F289", x"EE9A", x"ECBD", x"ED97", x"F11C", x"F6A6",
		x"FD44", x"03C6", x"091A", x"0C9A", x"0E81", x"0F37", x"0EE7", x"0D97",
		x"0B03", x"070D", x"01B5", x"FB60", x"F4FA", x"EF9A", x"EC90", x"EC91",
		x"EFCB", x"F53D", x"FB20", x"FFD5", x"023D", x"021D", x"0010", x"FC9D",
		x"F8BA", x"F4E9", x"F222", x"F0C2", x"F19A", x"F51D", x"FB14", x"029F",
		x"0A1D", x"0FD9", x"12D5", x"12F4", x"10DD", x"0DC1", x"0ABF", x"089C",
		x"073E", x"05EE", x"041A", x"012A", x"FD1E", x"F818", x"F306", x"EEF7",
		x"ECDF", x"ED78", x"F0C4", x"F60D", x"FC50", x"025E", x"0794", x"0B69",
		x"0E12", x"0FD1", x"110B", x"1239", x"1329", x"13FF", x"147A", x"14DB",
		x"1515", x"1521", x"14DD", x"1428", x"12D8", x"10A3", x"0D18", x"0802",
		x"0171", x"FA56", x"F3CD", x"EECF", x"EC62", x"ED31", x"F101", x"F741",
		x"FE9B", x"05DC", x"0C33", x"1122", x"13CF", x"13C4", x"10E6", x"0BAA",
		x"04DC", x"FD59", x"F617", x"F031", x"EC9F", x"EBB8", x"ED9C", x"F26D",
		x"F9D9", x"02CA", x"0B7F", x"119A", x"143C", x"143D", x"138F", x"1348",
		x"1359", x"12A7", x"0FE8", x"0AAA", x"031D", x"FAE9", x"F405", x"F092",
		x"F1D5", x"F734", x"FF5F", x"07B8", x"0E80", x"1265", x"13C3", x"13C6",
		x"1391", x"13C0", x"13C1", x"1274", x"0E85", x"07C6", x"FF1E", x"F679",
		x"EFD2", x"EC69", x"ECCB", x"F07C", x"F661", x"FD3F", x"041D", x"0A17",
		x"0ECD", x"1214", x"141E", x"1526", x"1562", x"151B", x"14A8", x"144E",
		x"13E3", x"132C", x"11E1", x"102A", x"0DFF", x"0B6F", x"0894", x"05A7",
		x"0302", x"00D1", x"FF19", x"FD83", x"FBE4", x"F9F8", x"F7AD", x"F506",
		x"F1CA", x"EE9E", x"EC1A", x"EB4B", x"ECF0", x"F0CA", x"F69F", x"FDAA",
		x"05A2", x"0CE4", x"11DE", x"131B", x"1025", x"09FD", x"024E", x"FAA5",
		x"F49B", x"F131", x"F10D", x"F47A", x"FAE6", x"02D1", x"0A79", x"1036",
		x"1367", x"1486", x"1499", x"1490", x"1492", x"13F2", x"118F", x"0C56",
		x"045F", x"FB52", x"F33C", x"EE1F", x"ED00", x"F009", x"F646", x"FE0D",
		x"0556", x"0AD1", x"0E03", x"0E98", x"0C6A", x"075F", x"0064", x"F8C2",
		x"F201", x"ED6A", x"EB9D", x"EC16", x"ED78", x"EE50", x"EDE2", x"ECC1",
		x"EBB4", x"EB58", x"EBF7", x"ED4E", x"EEFE", x"F09A", x"F1FC", x"F2F7",
		x"F403", x"F590", x"F822", x"FC0F", x"014D", x"074C", x"0D13", x"1175",
		x"136C", x"1270", x"0EC2", x"096E", x"03A1", x"FE2B", x"F9B8", x"F64A",
		x"F3F6", x"F26C", x"F12F", x"EFFA", x"EEAD", x"ED6D", x"EC63", x"EBB4",
		x"EB8A", x"EBEA", x"ECB3", x"ED61", x"ED4A", x"EC91", x"EC37", x"EDAC",
		x"F1F5", x"F8AC", x"00D7", x"08A1", x"0E6E", x"10D8", x"0F5A", x"09E2",
		x"01CA", x"F932", x"F20C", x"ED96", x"EBBD", x"EB6A", x"EB7C", x"EB72",
		x"EBA6", x"ED70", x"F1ED", x"F951", x"0242", x"0AB4", x"10B9", x"1328",
		x"11C1", x"0D10", x"0660", x"FF20", x"F88F", x"F386", x"F054", x"EEEA",
		x"EF32", x"F0BF", x"F337", x"F68B", x"FA30", x"FD3F", x"FF20", x"FF85",
		x"FE7D", x"FC82", x"F9D4", x"F6DD", x"F3DD", x"F182", x"EFBE", x"EED6",
		x"EEAC", x"EF24", x"F01F", x"F1B7", x"F420", x"F788", x"FC1D", x"0192",
		x"0771", x"0D01", x"1133", x"132F", x"12A4", x"0F6F", x"0A40", x"0413",
		x"FDBE", x"F84B", x"F42A", x"F181", x"EFBD", x"EE7F", x"ED9A", x"ED2E",
		x"ED72", x"EE62", x"EFD8", x"F1DC", x"F434", x"F69B", x"F8D5", x"FAA0",
		x"FBB0", x"FC4C", x"FC61", x"FBCE", x"FA54", x"F7EA", x"F4A7", x"F127",
		x"EE1B", x"EC62", x"ED14", x"F0A4", x"F6EB", x"FEB0", x"0671", x"0CA2",
		x"1070", x"116A", x"0F92", x"0B4F", x"04FE", x"FD6B", x"F5FA", x"F014",
		x"ECEA", x"ECB6", x"EED7", x"F1EC", x"F4D1", x"F71F", x"F8B9", x"F9AA",
		x"FA1F", x"FA6E", x"FAA0", x"FA90", x"FA12", x"F90A", x"F750", x"F4ED",
		x"F1E8", x"EEAD", x"EC5D", x"EC28", x"EEAD", x"F3F6", x"FB11", x"02C3",
		x"09C6", x"0F15", x"1228", x"1333", x"1270", x"108D", x"0DD0", x"0A9E",
		x"077A", x"0543", x"04CC", x"068C", x"0A94", x"0F60", x"12B0", x"12A1",
		x"0E9E", x"085F", x"0241", x"FE7A", x"FDB2", x"FF76", x"02FE", x"0754",
		x"0B55", x"0E97", x"103A", x"0F9A", x"0C4D", x"0653", x"FEAF", x"F6F1",
		x"F0A7", x"ECDE", x"EBBC", x"EC94", x"EE07", x"EF23", x"EF02", x"EDEC",
		x"EC65", x"EB1A", x"EAA4", x"EB12", x"EC38", x"EDA8", x"EF3F", x"F0C1",
		x"F264", x"F429", x"F63B", x"F87A", x"FB0B", x"FDDA", x"00CD", x"03B7",
		x"0677", x"08F5", x"0B28", x"0D44", x"0F1A", x"10A2", x"11E2", x"12EA",
		x"13E1", x"1497", x"14F9", x"14F4", x"148F", x"13E8", x"130B", x"1224",
		x"1142", x"1043", x"0EE7", x"0CB9", x"0936", x"0419", x"FD89", x"F661",
		x"F03E", x"EC99", x"EC49", x"EEC4", x"F288", x"F590", x"F684", x"F504",
		x"F1AC", x"EE43", x"ECE9", x"EF22", x"F4E6", x"FCE9", x"057A", x"0CDF",
		x"1215", x"1480", x"1415", x"10ED", x"0B9B", x"04D5", x"FD6B", x"F657",
		x"F0A7", x"ED1F", x"EC32", x"EDE3", x"F20F", x"F833", x"FFBA", x"0777",
		x"0E09", x"1247", x"130C", x"1099", x"0B86", x"059C", x"0082", x"FD53",
		x"FC9F", x"FE11", x"014C", x"0532", x"091C", x"0C37", x"0DF6", x"0DCE",
		x"0B60", x"0685", x"FFDE", x"F886", x"F208", x"EDD2", x"ECEC", x"EF6D",
		x"F4C5", x"FBC3", x"0341", x"0A34", x"0FA1", x"1327", x"1410", x"123B",
		x"0D92", x"06AD", x"FEC0", x"F72E", x"F11A", x"ED5E", x"EC27", x"ED28",
		x"EFBA", x"F329", x"F6E4", x"FA84", x"FDE8", x"0091", x"025C", x"0359",
		x"039C", x"0368", x"02FB", x"0249", x"0118", x"FF69", x"FCD8", x"F970",
		x"F51F", x"F0B7", x"EDA2", x"ECE6", x"EF52", x"F467", x"FB4A", x"0242",
		x"079D", x"0A0B", x"0950", x"05DD", x"0073", x"F9DD", x"F357", x"EE95",
		x"ED14", x"EFE9", x"F652", x"FEC5", x"074F", x"0E42", x"1295", x"1419",
		x"1390", x"11D7", x"105A", x"0FDF", x"10AD", x"1207", x"1375", x"146B",
		x"14D8", x"1537", x"1543", x"148F", x"126B", x"0E27", x"07AE", x"FF8F",
		x"F73A", x"F060", x"EC22", x"EA6F", x"EAAC", x"EC23", x"EE6F", x"F143",
		x"F420", x"F62A", x"F6CB", x"F59B", x"F2E7", x"EFA1", x"ED4B", x"ED44",
		x"F052", x"F5EC", x"FCED", x"03EA", x"09D4", x"0E53", x"1131", x"12E9",
		x"13BD", x"1422", x"1467", x"148B", x"1472", x"140B", x"1341", x"1232",
		x"10E5", x"0F49", x"0D1F", x"0A75", x"075A", x"03FE", x"00C8", x"FDCD",
		x"FB41", x"F8F6", x"F6B7", x"F48C", x"F2D3", x"F179", x"F027", x"EF02",
		x"EDE5", x"ECE9", x"EBED", x"EB1C", x"EAD6", x"EC15", x"EF87", x"F50A",
		x"FC26", x"03D2", x"0AFC", x"1062", x"1395", x"1449", x"1327", x"1117",
		x"0E8F", x"0C4D", x"0ABA", x"0A0B", x"0A51", x"0BB5", x"0E1E", x"10FC",
		x"1347", x"13B8", x"117D", x"0C60", x"04FD", x"FC96", x"F4C2", x"EF0C",
		x"EC10", x"EBC3", x"EDF8", x"F242", x"F87C", x"0015", x"07F5", x"0E73",
		x"1204", x"11F6", x"0EB3", x"0946", x"032E", x"FE5D", x"FC1B", x"FD5C",
		x"01A3", x"07BB", x"0DBA", x"11C4", x"12DB", x"10DD", x"0CB7", x"07B6",
		x"0346", x"003D", x"FE85", x"FDA4", x"FC95", x"FA9D", x"F75B", x"F312",
		x"EF18", x"ED0E", x"EDFF", x"F231", x"F87F", x"FF81", x"0514", x"07D3",
		x"06EC", x"027F", x"FBEC", x"F4D9", x"EF5E", x"ECC2", x"ED4D", x"F092",
		x"F527", x"F9B4", x"FCDD", x"FE91", x"FF49", x"0002", x"0218", x"05CE",
		x"0A88", x"0EE4", x"11A2", x"119E", x"0E72", x"08C7", x"0254", x"FD13",
		x"FAC2", x"FBF3", x"0037", x"0666", x"0CB7", x"1174", x"133B", x"11E5",
		x"0DF9", x"08BE", x"0339", x"FDFF", x"F9A0", x"F639", x"F3F9", x"F34E",
		x"F498", x"F811", x"FDA9", x"04B8", x"0BB4", x"10B1", x"12C9", x"1242",
		x"104F", x"0EE6", x"0F16", x"10C6", x"129D", x"1303", x"1044", x"0A4C",
		x"0282", x"FAB1", x"F434", x"EFA8", x"ECC8", x"EB53", x"EAF6", x"EB00",
		x"EB0F", x"EB16", x"EB88", x"ED62", x"F16E", x"F7BA", x"FF6A", x"0756",
		x"0E16", x"1289", x"14DF", x"1554", x"1542", x"14D5", x"1460", x"1376",
		x"120A", x"0FBA", x"0CA2", x"08E5", x"04EF", x"00FC", x"FD49", x"FA20",
		x"F7C1", x"F69E", x"F704", x"F961", x"FDCD", x"03F3", x"0AB8", x"1052",
		x"1318", x"12EA", x"109E", x"0D90", x"0B1A", x"09E7", x"0A97", x"0CAB",
		x"0F89", x"1238", x"1426", x"14F2", x"14F5", x"148C", x"141B", x"13CE",
		x"1361", x"128B", x"10F1", x"0E13", x"095B", x"02CA", x"FB08", x"F398",
		x"EE3F", x"EBF2", x"EC75", x"EE9B", x"F0E3", x"F267", x"F271", x"F136",
		x"EF4C", x"ED5B", x"EBC9", x"EAE9", x"EAA4", x"EAA2", x"EAB8", x"EAF4",
		x"EB1C", x"EB84", x"EC7C", x"EE57", x"F1BB", x"F6EB", x"FDB0", x"057C",
		x"0CC9", x"11CB", x"1387", x"1273", x"108D", x"0F79", x"101F", x"11CB",
		x"12F0", x"11E6", x"0DAE", x"06EA", x"FF59", x"F8EF", x"F4C6", x"F32F",
		x"F3AD", x"F5B7", x"F8D8", x"FCB9", x"0104", x"054A", x"095A", x"0CF9",
		x"0FEC", x"123B", x"13C2", x"1499", x"14F9", x"1503", x"148D", x"12E1",
		x"0F23", x"090C", x"015D", x"F961", x"F285", x"EDAA", x"EAFE", x"EA1F",
		x"EA52", x"EAC0", x"EB69", x"EC7B", x"EE48", x"F080", x"F24E", x"F2E9",
		x"F20B", x"F030", x"EE1B", x"EC83", x"EB81", x"EAC3", x"EA51", x"EA3F",
		x"EB76", x"EE65", x"F37A", x"FA9B", x"0280", x"09FC", x"0F9D", x"12F1",
		x"144D", x"146C", x"13E6", x"12F1", x"1133", x"0EC3", x"0C2F", x"0A24",
		x"0938", x"095F", x"0A6B", x"0C19", x"0E25", x"1036", x"1219", x"1393",
		x"149F", x"14EC", x"14AC", x"13FC", x"12DD", x"118E", x"1013", x"0EF8",
		x"0E79", x"0EAE", x"0F8F", x"10E6", x"1257", x"13A7", x"14A7", x"1540",
		x"156F", x"1570", x"1547", x"14FA", x"1498", x"13F8", x"133B", x"1232",
		x"10CE", x"0EBF", x"0BCC", x"0834", x"042F", x"004C", x"FCC3", x"FA3D",
		x"F94B", x"FA36", x"FD6A", x"0287", x"08A9", x"0E4D", x"1202", x"12CC",
		x"10B3", x"0C5E", x"0732", x"0240", x"FE23", x"FACD", x"F84A", x"F63A",
		x"F4C7", x"F37F", x"F248", x"F0FE", x"EFD0", x"EEAA", x"ED97", x"EC98",
		x"EB99", x"EB10", x"EBB3", x"EDA0", x"F153", x"F6B2", x"FD97", x"0515",
		x"0BF5", x"111A", x"13B1", x"140A", x"127E", x"0FE6", x"0CDF", x"09DD",
		x"07AB", x"06C5", x"0765", x"095C", x"0C39", x"0F7C", x"125C", x"13D8",
		x"12D4", x"0EC1", x"0804", x"FF8C", x"F70F", x"F074", x"ED34", x"EDF8",
		x"F212", x"F7C1", x"FD5E", x"00E9", x"0142", x"FE17", x"F857", x"F236",
		x"EDF1", x"ED00", x"EF4C", x"F2E8", x"F5A7", x"F5E4", x"F384", x"F009",
		x"EDBA", x"EE91", x"F2E8", x"F9C3", x"0132", x"0776", x"0BB4", x"0DE4",
		x"0EBA", x"0F00", x"0FA3", x"10EF", x"12D4", x"1427", x"13DA", x"10E3",
		x"0B2D", x"03BD", x"FBCE", x"F4D4", x"EFA2", x"ECA7", x"EB78", x"EB3A",
		x"EBC1", x"ED29", x"EF5D", x"F26B", x"F5FB", x"F98B", x"FCD2", x"FF76",
		x"0145", x"0282", x"038D", x"053C", x"0803", x"0BD3", x"0FEA", x"12B7",
		x"130F", x"104A", x"0AAB", x"037A", x"FC3B", x"F6C1", x"F430", x"F50A",
		x"F923", x"FF9B", x"06F0", x"0D67", x"11CA", x"1326", x"11AB", x"0E51",
		x"0A99", x"07EF", x"06B5", x"060E", x"04FA", x"029B", x"FEBD", x"F99E",
		x"F437", x"EFA1", x"ED7A", x"EE99", x"F2CB", x"F896", x"FDCF", x"0043",
		x"FEE5", x"FA42", x"F429", x"EF24", x"ED44", x"EEF5", x"F308", x"F78F",
		x"FA8E", x"FAF6", x"F8B3", x"F511", x"F138", x"EE52", x"EC8B", x"EBCF",
		x"ECBD", x"F048", x"F6AD", x"FEFB", x"0755", x"0E0E", x"125A", x"14AA",
		x"1581", x"1562", x"146A", x"11BC", x"0CC8", x"0580", x"FCD9", x"F4A4",
		x"EEA4", x"EB7F", x"EAA0", x"EB32", x"EC16", x"ED1C", x"EDEE", x"EE86",
		x"EEB8", x"EE6B", x"EDBF", x"ECF6", x"EC26", x"EB83", x"EB21", x"EB09",
		x"EB39", x"EB60", x"EB4D", x"EB00", x"EA9F", x"EA6F", x"EAAF", x"EB56",
		x"EC71", x"EE27", x"F0A4", x"F3C9", x"F788", x"FB41", x"FEBE", x"0177",
		x"02F1", x"027A", x"FFE8", x"FB45", x"F599", x"F03F", x"ED28", x"ED62",
		x"F076", x"F4DB", x"F8DB", x"FB28", x"FB5E", x"F9CB", x"F6D7", x"F37E",
		x"F095", x"EE96", x"ED66", x"ECB5", x"ECBC", x"ED47", x"EE4B", x"EFE9",
		x"F250", x"F5B0", x"FA24", x"FFCF", x"0606", x"0BF7", x"10AF", x"133C",
		x"1310", x"1058", x"0BB0", x"05E3", x"FFFD", x"FAD0", x"F6B2", x"F3A2",
		x"F16F", x"F01E", x"EF89", x"EF9E", x"F04D", x"F13B", x"F281", x"F413",
		x"F618", x"F873", x"FB47", x"FE4C", x"01A9", x"053F", x"092A", x"0D1D",
		x"1044", x"1259", x"136C", x"1359", x"11FB", x"0E82", x"08A1", x"00CA",
		x"F8A6", x"F1C5", x"ED1A", x"EAEC", x"EA85", x"EAC7", x"EB53", x"EC8A",
		x"EF8A", x"F507", x"FCDE", x"058E", x"0D05", x"120F", x"1453", x"14AC",
		x"13FB", x"12FB", x"11D1", x"1140", x"117A", x"127C", x"13B4", x"1409",
		x"1280", x"0E9F", x"0871", x"00EA", x"F94A", x"F306", x"EEB8", x"EC5D",
		x"EB76", x"EB65", x"EBBA", x"EC16", x"EC5C", x"EC4C", x"EC38", x"EC09",
		x"EBD5", x"EBC0", x"EC1E", x"ECC9", x"ED5C", x"ED51", x"ECA5", x"EBF0",
		x"EC01", x"EE03", x"F249", x"F8D7", x"0087", x"07FF", x"0DA2", x"10EE",
		x"1232", x"1235", x"113C", x"0F30", x"0C09", x"0791", x"0236", x"FC5D",
		x"F65F", x"F0DC", x"ED01", x"EB8E", x"ED03", x"F116", x"F6F2", x"FD6F",
		x"0384", x"085D", x"0BEA", x"0E4F", x"1005", x"1115", x"118E", x"1198",
		x"1125", x"1043", x"0ED4", x"0CEE", x"0A98", x"07FD", x"0586", x"036B",
		x"0219", x"019C", x"0201", x"035B", x"05B7", x"08EC", x"0C7E", x"0FD3",
		x"1270", x"13F5", x"1400", x"123B", x"0E2A", x"0808", x"0078", x"F8B6",
		x"F1F0", x"ED7A", x"EC30", x"EE49", x"F30F", x"F986", x"004F", x"069A",
		x"0BFE", x"1034", x"132B", x"14A7", x"1519", x"14BD", x"1433", x"13B8",
		x"137D", x"1370", x"13A5", x"13F1", x"143C", x"14A3", x"14D3", x"14DC",
		x"1437", x"1241", x"0E2F", x"078B", x"FF12", x"F683", x"EFD3", x"EC0E",
		x"EAE2", x"EAFB", x"EB4D", x"EBA5", x"ECEA", x"F003", x"F5A6", x"FD3D",
		x"0578", x"0C19", x"0F9E", x"0EFA", x"0A58", x"0323", x"FAF4", x"F3A8",
		x"EE95", x"EC19", x"EBCA", x"EC9D", x"ED35", x"ED06", x"EC2F", x"EB6A",
		x"EB4C", x"EBBE", x"EBE6", x"EBAE", x"EBB7", x"ED4A", x"F13F", x"F79D",
		x"FF6C", x"070F", x"0D56", x"1136", x"12C3", x"1273", x"10ED", x"0E92",
		x"0BC5", x"08D6", x"05FF", x"03D1", x"02BD", x"0302", x"0498", x"0701",
		x"09F5", x"0CAF", x"0F2B", x"114E", x"1315", x"1439", x"14C7", x"14C1",
		x"1450", x"139D", x"1313", x"12A4", x"126F", x"124C", x"126B", x"12EA",
		x"13BA", x"1497", x"1507", x"14AB", x"13AD", x"1257", x"10CB", x"0F51",
		x"0DAB", x"0C03", x"0A43", x"085D", x"05D5", x"029C", x"FECE", x"FA9B",
		x"F6BE", x"F379", x"F131", x"EFEE", x"EFAA", x"F0CD", x"F3D8", x"F919",
		x"002A", x"07A7", x"0E1F", x"1251", x"13E2", x"12E8", x"103F", x"0CE0",
		x"09F0", x"07E4", x"0658", x"04BC", x"0264", x"FF14", x"FAE2", x"F642",
		x"F1A1", x"EDF3", x"EC4E", x"EDB1", x"F240", x"F931", x"0138", x"08D1",
		x"0EDF", x"129F", x"1396", x"11CD", x"0DAE", x"080C", x"01BF", x"FB91",
		x"F63F", x"F234", x"EFA0", x"EE0B", x"ED1D", x"ECC1", x"ECF3", x"EE0A",
		x"F085", x"F4D4", x"FADF", x"0242", x"09BE", x"0FC3", x"12F1", x"126E",
		x"0ECA", x"0913", x"0260", x"FB94", x"F543", x"F01C", x"ECF0", x"EC70",
		x"EF07", x"F51C", x"FD89", x"069C", x"0E18", x"12CE", x"1504", x"15A4",
		x"1563", x"1496", x"1282", x"0E7D", x"0857", x"0094", x"F8B9", x"F230",
		x"EDF9", x"EBC5", x"EB17", x"EB58", x"EC20", x"ED9B", x"F02D", x"F45B",
		x"FA36", x"0159", x"08A9", x"0EF2", x"12C7", x"13A1", x"118C", x"0DD5",
		x"0A6D", x"08D9", x"09F2", x"0D35", x"10CF", x"12AF", x"113C", x"0C7A",
		x"0580", x"FE26", x"F7C9", x"F34C", x"F0BD", x"EFAA", x"EF3C", x"EECD",
		x"EE1E", x"ED23", x"EC28", x"EB7D", x"EB60", x"EC3E", x"EDB4", x"EF4E",
		x"F013", x"EFAE", x"EE3F", x"EC99", x"EBD8", x"ED25", x"F117", x"F75E",
		x"FED5", x"05EB", x"0BCE", x"0FEE", x"12B4", x"141F", x"14B2", x"14A3",
		x"1474", x"1491", x"1500", x"14F7", x"134E", x"0F1C", x"0870", x"0055",
		x"F843", x"F1A9", x"ED75", x"EC3E", x"EE15", x"F2ED", x"FA01", x"022A",
		x"0A31", x"105E", x"13DC", x"14F7", x"14C6", x"1469", x"1454", x"1410",
		x"1317", x"11A0", x"105C", x"1040", x"1144", x"12D9", x"139E", x"1229",
		x"0DC4", x"06EE", x"FF1E", x"F7E7", x"F237", x"EE43", x"EC07", x"EAF5",
		x"EA98", x"EA82", x"EA98", x"EB00", x"EBA1", x"EC84", x"EDA6", x"EF66",
		x"F1A1", x"F426", x"F648", x"F7BB", x"F827", x"F7C8", x"F684", x"F498",
		x"F281", x"F072", x"EED4", x"ED89", x"EC92", x"EBC1", x"EB4F", x"EB5F",
		x"EC16", x"ED49", x"EF33", x"F1FF", x"F5EC", x"FAEB", x"009B", x"06A0",
		x"0C52", x"1107", x"13C4", x"13D1", x"1080", x"0A41", x"0230", x"F9AE",
		x"F25E", x"ED74", x"EB96", x"ECC7", x"EFF8", x"F391", x"F66C", x"F7C3",
		x"F795", x"F625", x"F3A6", x"F0EB", x"EE72", x"EC97", x"EB66", x"EAC9",
		x"EA8D", x"EA87", x"EAB0", x"EB19", x"EBD4", x"ED6A", x"F067", x"F58E",
		x"FCE8", x"056A", x"0CF2", x"11AF", x"1356", x"12B9", x"11C7", x"1185",
		x"123E", x"133F", x"12D2", x"0FD8", x"09A6", x"01BD", x"FA1F", x"F4D8",
		x"F2B2", x"F373", x"F628", x"FA44", x"FEFB", x"0363", x"063F", x"0685",
		x"03A0", x"FDD1", x"F6A2", x"F08D", x"ED76", x"EE04", x"F0C8", x"F36C",
		x"F432", x"F2B8", x"EFEA", x"ED80", x"ED91", x"F13A", x"F778", x"FE80",
		x"041A", x"06F4", x"070A", x"04C2", x"00E2", x"FC5F", x"F838", x"F520",
		x"F369", x"F340", x"F46B", x"F6CF", x"FA04", x"FD68", x"00B6", x"0388",
		x"0577", x"0641", x"05F2", x"0475", x"024B", x"FFB5", x"FCC6", x"F9AD",
		x"F684", x"F391", x"F107", x"EEDB", x"ED1F", x"EBE0", x"EB4E", x"EB00",
		x"EAD8", x"EAA6", x"EA6F", x"EA73", x"EADA", x"EBE2", x"ED57", x"EF3F",
		x"F0E8", x"F1F6", x"F22F", x"F198", x"F053", x"EEB1", x"ED1B", x"EBE0",
		x"EB18", x"EAA9", x"EA85", x"EA7F", x"EA8C", x"EA8C", x"EAAB", x"EB2E",
		x"EC7F", x"EEE0", x"F287", x"F7A5", x"FE16", x"054A", x"0C08", x"1101",
		x"1369", x"1337", x"10C8", x"0D11", x"08D1", x"04E1", x"01AC", x"FF28",
		x"FD1B", x"FB47", x"F984", x"F7D7", x"F5D3", x"F3CA", x"F18F", x"EF8A",
		x"EDE4", x"EC95", x"EBB6", x"EB3F", x"EB2E", x"EB4A", x"EB96", x"EBCB",
		x"EBFD", x"ECA2", x"EE61", x"F1CC", x"F6EC", x"FDAA", x"052C", x"0C52",
		x"117C", x"13AD", x"1305", x"112A", x"0FEC", x"1022", x"11BA", x"136A",
		x"1384", x"10EF", x"0B31", x"0315", x"FA0D", x"F273", x"EDD3", x"ED1D",
		x"EFF2", x"F56B", x"FBE6", x"01E5", x"05F8", x"0707", x"0516", x"0090",
		x"FABC", x"F4B5", x"EFD0", x"ED86", x"EEFF", x"F42D", x"FC01", x"04A5",
		x"0C59", x"11C0", x"1418", x"13A4", x"1181", x"0F0F", x"0D7B", x"0D78",
		x"0EE2", x"10F9", x"12F5", x"1445", x"1507", x"1558", x"14E8", x"134D",
		x"0FFE", x"0AA7", x"0353", x"FAFA", x"F33F", x"EDA3", x"EAD8", x"EA5F",
		x"EB25", x"EC40", x"ED2E", x"EDE9", x"EEEE", x"F0AB", x"F3C9", x"F8A9",
		x"FEF5", x"062B", x"0CF3", x"11EF", x"13F8", x"1318", x"0FD8", x"0B5D",
		x"069B", x"0227", x"FE68", x"FB8A", x"F991", x"F82D", x"F752", x"F6FF",
		x"F737", x"F809", x"F95F", x"FB4C", x"FDF5", x"015A", x"0550", x"097B",
		x"0DB6", x"1136", x"134D", x"135D", x"108A", x"0B20", x"040F", x"FC4F",
		x"F524", x"EF85", x"EC6D", x"EC0D", x"EE54", x"F2E9", x"F907", x"0041",
		x"07B7", x"0E55", x"1299", x"13EA", x"1212", x"0DC7", x"07E5", x"0174",
		x"FB51", x"F5F2", x"F18E", x"EE2D", x"EBE9", x"EABF", x"EA4F", x"EA6A",
		x"EA9C", x"EBAE", x"EE6D", x"F3AC", x"FB27", x"037B", x"0B24", x"10E2",
		x"1467", x"15A8", x"14B2", x"1164", x"0BBD", x"0449", x"FC21", x"F4A3",
		x"EED3", x"EB8A", x"EAC9", x"EC15", x"EF36", x"F472", x"FBB3", x"043E",
		x"0C5A", x"11B5", x"1314", x"1053", x"0A5C", x"029F", x"FAB9", x"F408",
		x"EF17", x"EC33", x"EAE9", x"EA9D", x"EA99", x"EABD", x"EAF7", x"EBAD",
		x"ED1D", x"EF6C", x"F297", x"F63B", x"F9A9", x"FC96", x"FF2E", x"017C",
		x"0379", x"0504", x"05FC", x"06B0", x"0725", x"0710", x"0616", x"03FA",
		x"00D4", x"FCAB", x"F80E", x"F355", x"EF2E", x"EC92", x"EC1D", x"EE37",
		x"F28F", x"F8B5", x"FF88", x"061A", x"0BC6", x"0FE6", x"12A6", x"141C",
		x"14D6", x"152B", x"155F", x"154F", x"14E1", x"1332", x"0F70", x"0985",
		x"0218", x"FA62", x"F39E", x"EE9A", x"EBA4", x"EA79", x"EA61", x"EAD7",
		x"EB5D", x"EC4C", x"EE1A", x"F13E", x"F623", x"FCB0", x"0464", x"0BA5",
		x"10F5", x"1345", x"12D1", x"107D", x"0E19", x"0CEC", x"0DBD", x"1059",
		x"12C6", x"12F3", x"0FA6", x"0967", x"0198", x"FA32", x"F454", x"F075",
		x"EE54", x"ED50", x"ECCD", x"EC6C", x"EBEB", x"EB4B", x"EAB2", x"EA5C",
		x"EA54", x"EA98", x"EB2F", x"EC40", x"EDF3", x"F0AA", x"F4A0", x"FA22",
		x"00EE", x"081D", x"0E38", x"1227", x"13A3", x"129D", x"0F61", x"0ADD",
		x"05E7", x"0129", x"FD3D", x"FA39", x"F84C", x"F7DB", x"F957", x"FD35",
		x"0325", x"0A06", x"0FAC", x"127B", x"11E0", x"0EF9", x"0C3C", x"0B5E",
		x"0D1F", x"1046", x"1283", x"11BB", x"0D4E", x"0683", x"FFFD", x"FC74",
		x"FD4B", x"023F", x"0925", x"0F33", x"120A", x"1142", x"0E1A", x"0B36",
		x"0A82", x"0C6E", x"0FC2", x"1292", x"128B", x"0ED4", x"0841", x"0088",
		x"F994", x"F47E", x"F13D", x"EF4D", x"EE14", x"ED1C", x"EC69", x"EBCD",
		x"EB37", x"EAB7", x"EA81", x"EAEB", x"EC28", x"EDB6", x"EF10", x"EFED",
		x"F04E", x"F042", x"EFED", x"EF11", x"EDF6", x"ECAC", x"EB9E", x"EAF8",
		x"EABB", x"EB0E", x"EBAF", x"ECA6", x"EDA1", x"EE77", x"EF70", x"F11B",
		x"F439", x"F8F2", x"FF6A", x"06CA", x"0D8F", x"1204", x"1314", x"1115",
		x"0DC5", x"0B50", x"0B37", x"0D58", x"1096", x"12D9", x"1266", x"0EB4",
		x"08B2", x"0213", x"FCAB", x"F965", x"F886", x"F9CB", x"FCBC", x"00EA",
		x"05A6", x"0A4B", x"0E8F", x"11E4", x"13E5", x"13F0", x"1177", x"0C90",
		x"05B9", x"FDE5", x"F639", x"F031", x"ECEB", x"ED56", x"F12F", x"F770",
		x"FE7F", x"04FC", x"09CD", x"0C8B", x"0D47", x"0C25", x"09C8", x"0686",
		x"02C7", x"FEFA", x"FC13", x"FAAE", x"FB37", x"FD84", x"0102", x"04FE",
		x"08B5", x"0B9D", x"0D2D", x"0D4A", x"0B79", x"07A7", x"01E3", x"FAEB",
		x"F412", x"EED2", x"EC60", x"ED80", x"F246", x"F9BC", x"026E", x"0A74",
		x"1069", x"13AE", x"1468", x"1388", x"11ED", x"10BE", x"108E", x"112B",
		x"1251", x"134E", x"13C8", x"1416", x"1440", x"1497", x"14C5", x"14B4",
		x"1434", x"134B", x"1238", x"111D", x"1048", x"1000", x"1097", x"11F6",
		x"13B9", x"14FD", x"1560", x"1519", x"14D0", x"14CD", x"14A3", x"1310",
		x"0F33", x"08C7", x"00C3", x"F885", x"F1AA", x"ED52", x"EB94", x"EB9C",
		x"ECE8", x"EEE1", x"F175", x"F47B", x"F782", x"F9D7", x"FAD9", x"FA6C",
		x"F888", x"F5B9", x"F2A1", x"EFEE", x"EDCA", x"ECAA", x"EC5E", x"ECA0",
		x"ED35", x"EE0F", x"EF2E", x"F0F1", x"F38E", x"F6B5", x"F9EE", x"FD56",
		x"00C2", x"0430", x"0762", x"0A09", x"0C0B", x"0D7B", x"0E56", x"0EB1",
		x"0E78", x"0DB7", x"0C25", x"09BF", x"06D1", x"03BC", x"0097", x"FD4D",
		x"F9DC", x"F693", x"F3CA", x"F193", x"EFD3", x"EE8B", x"ED95", x"ED19",
		x"ECEF", x"ED08", x"ED80", x"EE58", x"EFE3", x"F205", x"F530", x"F97A",
		x"FF07", x"05A7", x"0C16", x"110A", x"136F", x"130C", x"100C", x"0B7A",
		x"0622", x"0120", x"FD2A", x"FA5C", x"F867", x"F6AF", x"F4CF", x"F291",
		x"F008", x"EDA8", x"EC0E", x"EC65", x"EF6C", x"F54E", x"FD0F", x"04FC",
		x"0B80", x"0FEC", x"127A", x"13C6", x"1460", x"1496", x"14A6", x"14BC",
		x"146F", x"12CF", x"0F02", x"08D0", x"00A1", x"F84D", x"F157", x"ECDE",
		x"EB03", x"EA83", x"EAC7", x"EB2A", x"EC54", x"EF43", x"F4DC", x"FCD5",
		x"05C7", x"0DA9", x"12AB", x"1409", x"120A", x"0D64", x"070D", x"FFED",
		x"F8FC", x"F2CF", x"EE55", x"EC1B", x"ECBB", x"F00E", x"F59E", x"FC7C",
		x"03D9", x"0AB4", x"1025", x"134D", x"13A5", x"10EA", x"0BA9", x"04D1",
		x"FD68", x"F671", x"F0E5", x"ED0F", x"EAE8", x"EA69", x"EAE1", x"EBF6",
		x"ED00", x"ED93", x"ED8B", x"ECDE", x"EBE7", x"EB7E", x"EC7F", x"EFB6",
		x"F5B3", x"FD9D", x"0635", x"0D84", x"1243", x"13EF", x"12B9", x"0EF6",
		x"091C", x"01E1", x"FA54", x"F396", x"EE9D", x"EC0E", x"EC41", x"EF00",
		x"F3D4", x"FA25", x"0145", x"0891", x"0ECB", x"12DB", x"1399", x"10AE",
		x"0ACC", x"0359", x"FC13", x"F62C", x"F228", x"EFCA", x"EEAD", x"EE90",
		x"EF2D", x"F097", x"F322", x"F72C", x"FCB5", x"034A", x"0A26", x"0FB4",
		x"12D2", x"12B2", x"0FB0", x"0B36", x"06F3", x"048B", x"04C2", x"078E",
		x"0BE6", x"102A", x"127D", x"1156", x"0C89", x"0500", x"FC54", x"F462",
		x"EEB2", x"EBDE", x"EBDD", x"EE48", x"F28D", x"F7EB", x"FDCC", x"0376",
		x"08B1", x"0CF0", x"1023", x"11EC", x"128B", x"1212", x"104A", x"0D2F",
		x"0837", x"01CF", x"FA8F", x"F397", x"EE46", x"EB93", x"EBB6", x"EE43",
		x"F24E", x"F6B4", x"FA9C", x"FD79", x"FF3A", x"FF6A", x"FE17", x"FB76",
		x"F7C0", x"F370", x"EF7E", x"ECE6", x"ECC2", x"EFB8", x"F59B", x"FDA5",
		x"062D", x"0D96", x"1267", x"13B4", x"11BE", x"0DCC", x"095E", x"0584",
		x"02C8", x"0128", x"00D4", x"01E9", x"0445", x"0794", x"0B69", x"0F49",
		x"1257", x"13C2", x"12E6", x"0F5D", x"097B", x"0243", x"FAE4", x"F462",
		x"EFAA", x"ECCA", x"EB6E", x"EB03", x"EAF2", x"EAE7", x"EAF7", x"EB48",
		x"EC7C", x"EF9D", x"F534", x"FCEE", x"0542", x"0C87", x"1180", x"13F6",
		x"1486", x"140F", x"13AA", x"13C1", x"1440", x"1474", x"140D", x"137C",
		x"1329", x"1365", x"1407", x"145E", x"135E", x"1022", x"0A30", x"023D",
		x"F9A6", x"F234", x"ED47", x"EB6E", x"ECB8", x"F0A4", x"F674", x"FD68",
		x"04D4", x"0BA1", x"10CA", x"136A", x"12DC", x"0F47", x"0973", x"0257",
		x"FB20", x"F4D1", x"F020", x"ED03", x"EB67", x"EABC", x"EA9D", x"EAEA",
		x"EB5C", x"EBC7", x"EC32", x"ECE6", x"EDCB", x"EEC5", x"EFCD", x"F106",
		x"F2E3", x"F5F3", x"FA94", x"009A", x"0763", x"0DAE", x"11FC", x"134B",
		x"1190", x"0DDE", x"09D5", x"0756", x"0752", x"09FB", x"0E13", x"11B4",
		x"132D", x"1124", x"0B94", x"037F", x"FA71", x"F2A6", x"EDCD", x"ECD5",
		x"EF5B", x"F41C", x"F91D", x"FC93", x"FD1D", x"FA3E", x"F50F", x"EFDD",
		x"ECFA", x"EDCD", x"F1B2", x"F684", x"F9B1", x"F991", x"F664", x"F1B5",
		x"EE69", x"EE76", x"F25D", x"F82E", x"FDB9", x"0112", x"0192", x"FF92",
		x"FBE5", x"F7A6", x"F3C8", x"F0F6", x"EFE4", x"F0F7", x"F4B3", x"FAD1",
		x"022E", x"0999", x"0F8F", x"12F1", x"1373", x"11A8", x"0E7D", x"0B0F",
		x"0808", x"0587", x"036B", x"017E", x"FFD3", x"FE1A", x"FC2E", x"F9FE",
		x"F793", x"F543", x"F327", x"F14F", x"EF75", x"EDC9", x"EC92", x"EBDD",
		x"EB7B", x"EB6E", x"EB9C", x"EC0E", x"ECC3", x"ED77", x"EE23", x"EE5E",
		x"EE21", x"ED69", x"EC72", x"EB85", x"EB06", x"EB46", x"EC63", x"EED3",
		x"F2AE", x"F832", x"FEFE", x"0630", x"0C9E", x"113E", x"1343", x"11D8",
		x"0CD9", x"0505", x"FBFE", x"F40A", x"EE8C", x"EBA3", x"EA93", x"EA62",
		x"EAA7", x"EBBF", x"EE94", x"F3A2", x"FAF6", x"0364", x"0B44", x"10FD",
		x"13F6", x"14E3", x"14BC", x"1494", x"1485", x"1453", x"13C6", x"1239",
		x"0EBE", x"08B9", x"009D", x"F7E4", x"F102", x"ED31", x"EC33", x"EC9E",
		x"ED07", x"ECE5", x"ECA6", x"ED62", x"F047", x"F59B", x"FCDF", x"047D",
		x"0ABD", x"0E87", x"101F", x"0FFB", x"0EFF", x"0D21", x"0A2B", x"05CD",
		x"0021", x"F998", x"F35B", x"EEAC", x"ECB6", x"EE2D", x"F29A", x"F844",
		x"FD48", x"FFB1", x"FED0", x"FB05", x"F587", x"F069", x"ED7C", x"EDCA",
		x"F133", x"F6A1", x"FCBE", x"0279", x"0716", x"0A6A", x"0C94", x"0DDF",
		x"0E75", x"0EA0", x"0E01", x"0C95", x"0A38", x"06DF", x"0310", x"FFA3",
		x"FD55", x"FC84", x"FDB9", x"00F1", x"05F8", x"0BA9", x"1096", x"1317",
		x"128D", x"0F40", x"09F1", x"03C0", x"FD9B", x"F870", x"F48A", x"F205",
		x"F0B2", x"F059", x"F151", x"F3BC", x"F83E", x"FEAD", x"0629", x"0D2D",
		x"11D6", x"13A6", x"1317", x"114A", x"0FD4", x"0F9F", x"109A", x"1245",
		x"13C1", x"14B7", x"14F0", x"150E", x"1515", x"1517", x"150E", x"145A",
		x"1312", x"1170", x"1037", x"100C", x"1100", x"1284", x"13A2", x"12EB",
		x"0F76", x"0932", x"014C", x"F995", x"F343", x"EF09", x"EC78", x"EB58",
		x"EB0D", x"EAEC", x"EAFA", x"EB1C", x"EB75", x"EBE3", x"EC99", x"ED95",
		x"EF0C", x"F0D4", x"F2DE", x"F4DF", x"F715", x"F9B4", x"FCD0", x"0044",
		x"03F5", x"0786", x"0A78", x"0C9C", x"0DAC", x"0DAE", x"0C97", x"0A59",
		x"0710", x"0371", x"FFF4", x"FD6D", x"FC04", x"FC37", x"FE3D", x"0238",
		x"0774", x"0CE8", x"1171", x"1367", x"11FF", x"0CEA", x"051D", x"FC41",
		x"F43E", x"EED9", x"EC83", x"ED34", x"EFB4", x"F28E", x"F40D", x"F36B",
		x"F103", x"EE15", x"EC93", x"EE05", x"F2AF", x"F9C1", x"015C", x"0805",
		x"0CC3", x"0FBB", x"1149", x"1215", x"1297", x"132D", x"13E5", x"1478",
		x"14CF", x"1473", x"1357", x"11A8", x"0FB1", x"0E3A", x"0DF3", x"0F1D",
		x"113E", x"1320", x"132D", x"1082", x"0B27", x"046E", x"FD70", x"F793",
		x"F3D0", x"F22D", x"F244", x"F35C", x"F572", x"F8BE", x"FD6C", x"034D",
		x"0978", x"0EC9", x"1220", x"1278", x"0FC4", x"0AAB", x"0484", x"FF3D",
		x"FCC5", x"FDF8", x"029A", x"0926", x"0F23", x"1278", x"1270", x"0FD6",
		x"0C35", x"093B", x"0807", x"08DA", x"0B49", x"0E71", x"114F", x"1351",
		x"145A", x"14E4", x"1503", x"14BF", x"1432", x"133D", x"11D2", x"0F91",
		x"0C19", x"0764", x"017A", x"FAFE", x"F484", x"EF3E", x"EC30", x"EC12",
		x"EEBA", x"F36F", x"F8D5", x"FE09", x"0262", x"0592", x"07F4", x"09B9",
		x"0B06", x"0BA3", x"0B96", x"0A8D", x"089D", x"05BF", x"0255", x"FECF",
		x"FBBD", x"F989", x"F872", x"F8CB", x"FACD", x"FE6F", x"02C5", x"0704",
		x"0A53", x"0BF4", x"0B85", x"0866", x"02A3", x"FB0B", x"F3AB", x"EE89",
		x"EC88", x"ED2D", x"EEAF", x"EF8A", x"EEF7", x"ED6F", x"EC83", x"EDDE",
		x"F286", x"F9AE", x"01C1", x"08F3", x"0E5B", x"11CD", x"13E1", x"14CD",
		x"1522", x"1563", x"159A", x"15B6", x"15B4", x"1585", x"154C", x"14D0",
		x"1404", x"129B", x"1097", x"0E47", x"0BAE", x"08D3", x"05AB", x"0219",
		x"FE77", x"FB54", x"F91D", x"F7F7", x"F7E7", x"F8E9", x"FB2B", x"FE81",
		x"025A", x"0614", x"0907", x"0ABB", x"0AA5", x"0814", x"02CD", x"FB96",
		x"F449", x"EEDF", x"EC92", x"ED75", x"F01E", x"F28D", x"F382", x"F2A2",
		x"F0AA", x"EE5E", x"EC79", x"EB49", x"EA94", x"EA64", x"EB14", x"ED8D",
		x"F269", x"F974", x"0175", x"093E", x"0F94", x"1385", x"151C", x"14EA",
		x"13D3", x"129A", x"1166", x"1031", x"0ECB", x"0D3A", x"0B2A", x"08B5",
		x"05A6", x"0228", x"FEAC", x"FB80", x"F908", x"F782", x"F6EF", x"F743",
		x"F88A", x"FAA7", x"FD55", x"007F", x"03E2", x"0734", x"0A0E", x"0C21",
		x"0D93", x"0EDF", x"1049", x"11DC", x"1325", x"1444", x"14F0", x"14B5",
		x"1317", x"0F99", x"0A37", x"0369", x"FC18", x"F4FE", x"EF72", x"EC9A",
		x"ED77", x"F206", x"F939", x"014C", x"08AE", x"0E6F", x"1213", x"1428",
		x"1511", x"1550", x"156C", x"1550", x"1487", x"12EB", x"0FF9", x"0BDC",
		x"06AE", x"00AA", x"FA72", x"F47E", x"EF94", x"EC78", x"EC15", x"EEE8",
		x"F4C5", x"FCC3", x"0567", x"0CE1", x"11A6", x"1337", x"1206", x"0FB9",
		x"0E25", x"0E5D", x"104D", x"1262", x"12AE", x"1019", x"0A46", x"0322",
		x"FC6E", x"F80B", x"F6A6", x"F7F5", x"FB13", x"FF57", x"03B2", x"0753",
		x"0975", x"0972", x"0718", x"026E", x"FC2C", x"F56E", x"EFCE", x"ECAC",
		x"ED22", x"F14E", x"F845", x"00C1", x"091B", x"0FC4", x"136C", x"144D",
		x"130B", x"10B1", x"0EA7", x"0D6E", x"0D5E", x"0E27", x"0FA0", x"117D",
		x"1332", x"1472", x"14B4", x"142E", x"1311", x"1196", x"1001", x"0E76",
		x"0D49", x"0C71", x"0BB1", x"0B12", x"0AD8", x"0B38", x"0C65", x"0E38",
		x"107D", x"12C1", x"1485", x"14CB", x"12F3", x"0E58", x"0755", x"FF1B",
		x"F727", x"F0F2", x"ED04", x"EB13", x"EA96", x"EB3F", x"EC9A", x"EEB3",
		x"F143", x"F3D7", x"F57B", x"F578", x"F375", x"F067", x"EDB4", x"ECEE",
		x"EEFD", x"F3F8", x"FA7D", x"00F6", x"05A7", x"0800", x"086C", x"0748",
		x"051A", x"01BF", x"FD66", x"F83A", x"F322", x"EEDA", x"EC7D", x"ECBA",
		x"EFC7", x"F53E", x"FC24", x"0317", x"0854", x"0B72", x"0C54", x"0B84",
		x"0972", x"0648", x"0277", x"FE48", x"FA59", x"F6B9", x"F3CE", x"F16D",
		x"EFAF", x"EE66", x"ED6C", x"EC9B", x"EBCD", x"EAFE", x"EA6A", x"EA5A",
		x"EACD", x"EB66", x"EC28", x"ED36", x"EEEC", x"F1E3", x"F64F", x"FC55",
		x"0380", x"0ABD", x"107B", x"139D", x"139B", x"1129", x"0D62", x"09AD",
		x"06AF", x"04EA", x"03E8", x"02F9", x"014F", x"FDF9", x"F924", x"F3AF",
		x"EF47", x"ED2C", x"EE3E", x"F23C", x"F7F9", x"FD90", x"0129", x"01D6",
		x"FF69", x"FABC", x"F50A", x"EFD9", x"ED1C", x"EDF5", x"F2B5", x"FA81",
		x"0379", x"0B98", x"1128", x"138C", x"12F6", x"1071", x"0DB0", x"0C11",
		x"0C69", x"0E9F", x"1185", x"1337", x"124D", x"0E2A", x"0723", x"FE98",
		x"F64A", x"EFB0", x"EC0F", x"EBB4", x"EE4E", x"F2FA", x"F8A7", x"FEC3",
		x"04B5", x"09FD", x"0E2E", x"1146", x"134A", x"146B", x"14E7", x"14DD",
		x"142E", x"1219", x"0E08", x"07D1", x"001A", x"F83C", x"F18E", x"ED0D",
		x"EB13", x"EB3E", x"ECBF", x"EEA9", x"F070", x"F1E9", x"F35B", x"F52F",
		x"F7DA", x"FBB4", x"00CE", x"06DD", x"0CC8", x"117C", x"139D", x"1274",
		x"0E2C", x"0729", x"FEC7", x"F6B5", x"F059", x"EC9A", x"EBE7", x"EDCD",
		x"F128", x"F4CE", x"F7CA", x"F953", x"F95F", x"F7E0", x"F527", x"F1D1",
		x"EE8F", x"EC2F", x"EB43", x"EC0D", x"EE7D", x"F2D1", x"F8BA", x"0014",
		x"07B8", x"0E49", x"128C", x"13AE", x"1198", x"0D20", x"0721", x"005E",
		x"F99E", x"F390", x"EEF2", x"ECCD", x"EE20", x"F2E8", x"FA42", x"029E",
		x"0A22", x"0FC3", x"131F", x"145A", x"141A", x"12C2", x"109C", x"0DEB",
		x"0B0B", x"08A5", x"078B", x"0822", x"0A93", x"0E0C", x"1176", x"1384",
		x"12FC", x"0F5E", x"08D8", x"0061", x"F7B4", x"F0C6", x"ED01", x"ED19",
		x"F07B", x"F5B6", x"FB06", x"FEC3", x"FFBF", x"FDAC", x"F91D", x"F382",
		x"EED5", x"ECBA", x"EDEE", x"F21D", x"F80B", x"FE7C", x"03E5", x"07D8",
		x"0A56", x"0BC8", x"0CCF", x"0D72", x"0DAF", x"0D7C", x"0CFF", x"0C89",
		x"0C0E", x"0AEA", x"089E", x"04DF", x"FF8A", x"F95F", x"F36E", x"EEC9",
		x"ECBE", x"ED9E", x"F12F", x"F658", x"FBA4", x"FFD7", x"0274", x"03B0",
		x"0370", x"01BF", x"FEC9", x"FAD5", x"F65D", x"F1E8", x"EE33", x"EC3F",
		x"ED2B", x"F123", x"F77A", x"FEC9", x"05A3", x"0AF8", x"0E25", x"0EE6",
		x"0D95", x"0A99", x"06C6", x"02E6", x"FF86", x"FDA9", x"FE2B", x"0166",
		x"06D7", x"0CE5", x"115E", x"12DD", x"111D", x"0D42", x"0902", x"05A1",
		x"03E4", x"0405", x"05D2", x"08B5", x"0C30", x"0F83", x"1242", x"1402",
		x"1407", x"11E7", x"0D5B", x"06F5", x"FF81", x"F847", x"F24B", x"EDDB",
		x"EB58", x"EA72", x"EAAD", x"EB5D", x"EC0B", x"EC9B", x"ED2A", x"EDF5",
		x"EF53", x"F163", x"F3E7", x"F6AB", x"F999", x"FC75", x"FF33", x"01B9",
		x"0409", x"0602", x"07BF", x"0991", x"0B74", x"0DA5", x"0FD4", x"1214",
		x"13EE", x"14DB", x"1423", x"114F", x"0C22", x"0511", x"FD27", x"F578",
		x"EF86", x"EC38", x"EC03", x"EEAB", x"F383", x"F9A1", x"005C", x"0751",
		x"0D9E", x"11EB", x"12F0", x"0FE6", x"0987", x"018D", x"F9DC", x"F3B4",
		x"EFE7", x"EE9C", x"EFAB", x"F2D0", x"F7D4", x"FE4C", x"05C0", x"0CED",
		x"11EF", x"130D", x"0F9E", x"0847", x"FF0E", x"F673", x"F02B", x"EC93",
		x"EB11", x"EA9A", x"EA8B", x"EB28", x"ED14", x"F13C", x"F7B0", x"FF92",
		x"075E", x"0DA0", x"1109", x"1105", x"0DD8", x"0801", x"0076", x"F869",
		x"F160", x"ECD3", x"EBA0", x"ED52", x"F01B", x"F2A4", x"F407", x"F4D1",
		x"F5C1", x"F7E4", x"FB7B", x"0079", x"0673", x"0C80", x"113C", x"1371",
		x"128D", x"0EEB", x"09CB", x"0452", x"FF85", x"FB7F", x"F823", x"F57C",
		x"F358", x"F1A7", x"F044", x"EEFD", x"EDCE", x"ECF3", x"EC47", x"EBCA",
		x"EB6B", x"EB3D", x"EB6F", x"EC68", x"EF15", x"F3E7", x"FAF4", x"0323",
		x"0AD5", x"1084", x"13B4", x"14E7", x"151A", x"1509", x"14D6", x"13A6",
		x"1023", x"09A9", x"0119", x"F815", x"F0F6", x"ECD7", x"EC30", x"EE54",
		x"F2A8", x"F883", x"FF0E", x"0604", x"0C8B", x"115D", x"130B", x"1083",
		x"0A7B", x"0299", x"FAD8", x"F48C", x"F088", x"EF41", x"F10C", x"F5BD",
		x"FC9A", x"0474", x"0BAA", x"111B", x"1434", x"1509", x"14AB", x"1421",
		x"140F", x"146D", x"14AD", x"1448", x"138D", x"1315", x"1360", x"1415",
		x"1447", x"12B6", x"0E73", x"075C", x"FEB1", x"F622", x"EFBE", x"EC9D",
		x"EC9F", x"EF89", x"F4B4", x"FBA8", x"0305", x"0993", x"0E99", x"11EB",
		x"13DB", x"14BC", x"1518", x"152A", x"14E8", x"1472", x"137C", x"1228",
		x"1093", x"0E5A", x"0BAB", x"08D9", x"0644", x"0408", x"028A", x"01A2",
		x"0175", x"0222", x"037B", x"0530", x"0720", x"09D3", x"0D0D", x"1080",
		x"12E5", x"1316", x"105B", x"0AD4", x"0386", x"FBBC", x"F51B", x"F0C0",
		x"EFCE", x"F2F0", x"F9B4", x"0235", x"0A1F", x"0FD2", x"1317", x"145B",
		x"149A", x"1462", x"13C0", x"121A", x"0E36", x"07CF", x"FF95", x"F7A2",
		x"F188", x"EE21", x"ED1F", x"ED93", x"EEE6", x"F116", x"F428", x"F837",
		x"FD52", x"036D", x"09C7", x"0F45", x"1294", x"12EE", x"107D", x"0BD6",
		x"06A4", x"0252", x"0018", x"0031", x"0244", x"0575", x"0913", x"0C73",
		x"0F0A", x"109D", x"1121", x"10BC", x"0F81", x"0DC5", x"0B7A", x"08B4",
		x"059F", x"0214", x"FE22", x"FA19", x"F63C", x"F2E0", x"F056", x"EEA1",
		x"ED7E", x"ED10", x"EDB1", x"F030", x"F4E1", x"FB99", x"0336", x"0A94",
		x"106D", x"13B3", x"1424", x"1275", x"0FB1", x"0D3A", x"0B52", x"09F1",
		x"08B7", x"0773", x"05AD", x"02F6", x"FF4A", x"FB04", x"F6DB", x"F347",
		x"F0AE", x"EF5B", x"EF64", x"F0F4", x"F429", x"F91D", x"FFA7", x"06DD",
		x"0D43", x"11AB", x"1377", x"129D", x"0FA5", x"0B5E", x"06C7", x"02AD",
		x"FFBB", x"FE4A", x"FE36", x"FF89", x"022E", x"05FA", x"0A7D", x"0F06",
		x"1277", x"13BE", x"11B9", x"0C61", x"0473", x"FB99", x"F3D4", x"EEAE",
		x"ECA7", x"EDBF", x"F10C", x"F50A", x"F879", x"FA5A", x"FA2B", x"F840",
		x"F54E", x"F22E", x"EFBF", x"EE24", x"ED67", x"EDEC", x"F043", x"F4E3",
		x"FBB7", x"03BF", x"0B79", x"114A", x"146C", x"149C", x"12BF", x"1058",
		x"0E84", x"0D76", x"0CB2", x"0B72", x"0910", x"051C", x"FF8E", x"F8D4",
		x"F257", x"EDC3", x"EC6F", x"EE7D", x"F264", x"F678", x"F94E", x"FA64",
		x"F9D4", x"F7E0", x"F530", x"F24E", x"EFDD", x"EDFE", x"ECCB", x"EC55",
		x"EC56", x"ECF4", x"EE3A", x"F03B", x"F317", x"F6EA", x"FBC5", x"0153",
		x"072A", x"0C8B", x"10E4", x"137A", x"1379", x"109E", x"0AEB", x"032F",
		x"FADD", x"F363", x"EE2B", x"EBC6", x"EC6F", x"EF77", x"F3DC", x"F8E1",
		x"FDB8", x"0215", x"0576", x"07D3", x"0971", x"0AD8", x"0C51", x"0E0E",
		x"0FEA", x"11C7", x"1370", x"147D", x"14B8", x"1481", x"145A", x"14CB",
		x"153E", x"1470", x"113A", x"0B30", x"034D", x"FB1F", x"F403", x"EEBD",
		x"EC3D", x"ED59", x"F228", x"F9CB", x"0259", x"0A0D", x"1012", x"1412",
		x"161E", x"1627", x"1435", x"1082", x"0AFF", x"03A3", x"FB54", x"F361",
		x"EDC4", x"EBAD", x"ED66", x"F26C", x"F9C2", x"0241", x"0A66", x"10BE",
		x"147E", x"15D3", x"15AC", x"1515", x"14A0", x"1437", x"1387", x"126D",
		x"10F5", x"100A", x"0FF2", x"10AF", x"11D2", x"130D", x"1409", x"1496",
		x"14D7", x"14DD", x"14E4", x"1502", x"1528", x"150D", x"149F", x"13BE",
		x"1264", x"10DF", x"0F1C", x"0CF5", x"0A63", x"07F0", x"059F", x"038B",
		x"0165", x"FECC", x"FBF2", x"F8D4", x"F5D6", x"F2F7", x"F061", x"EE59",
		x"ECF5", x"EC2B", x"EBD0", x"EBE2", x"EC42", x"ED11", x"EE52", x"F037",
		x"F290", x"F4D5", x"F6AE", x"F7DE", x"F853", x"F7D3", x"F6A3", x"F4C6",
		x"F29F", x"F030", x"EDCD", x"EC0B", x"EB6D", x"ECB6", x"EFFC", x"F536",
		x"FBFE", x"0396", x"0ABC", x"103D", x"1321", x"12A6", x"0F02", x"08DC",
		x"0129", x"F993", x"F33E", x"EEDC", x"EC32", x"EB16", x"EAE4", x"EB4D",
		x"EC49", x"ED84", x"EED9", x"F030", x"F163", x"F2B3", x"F43D", x"F5E2",
		x"F76F", x"F936", x"FB8F", x"FF07", x"03A7", x"090B", x"0E26", x"11BD",
		x"12A2", x"102C", x"0AEB", x"0470", x"FEF7", x"FC79", x"FE17", x"0352",
		x"0A3A", x"0FF4", x"126C", x"1174", x"0E7B", x"0BDF", x"0B85", x"0D83",
		x"1061", x"11CB", x"0FCE", x"0A5F", x"032F", x"FD41", x"FB4E", x"FE35",
		x"04C3", x"0C29", x"1171", x"1306", x"1136", x"0E07", x"0BE4", x"0C51",
		x"0EDF", x"11BD", x"1281", x"0FD5", x"0A0E", x"032F", x"FD14", x"F95C",
		x"F857", x"F9D6", x"FD05", x"0101", x"04E0", x"0852", x"0AC7", x"0C0A",
		x"0BFB", x"0A9F", x"0842", x"0512", x"0180", x"FE05", x"FAD1", x"F814",
		x"F5AD", x"F389", x"F193", x"EFBF", x"EE39", x"ECF0", x"EBEC", x"EB34",
		x"EAB7", x"EAB3", x"EB21", x"EBF6", x"ED0A", x"EE3F", x"EF95", x"F13E",
		x"F36A", x"F65C", x"FA00", x"FDE7", x"0166", x"0437", x"063E", x"076D",
		x"07A8", x"0693", x"043F", x"0102", x"FD6D", x"FA1E", x"F765", x"F5C2",
		x"F58E", x"F771", x"FB8E", x"01A2", x"0888", x"0E91", x"1242", x"12A4",
		x"0FA0", x"09BE", x"026C", x"FAF0", x"F444", x"EF5E", x"EC96", x"EC73",
		x"EEE9", x"F3E8", x"FACC", x"029B", x"0A0C", x"0FD0", x"1319", x"13BA",
		x"1225", x"0F13", x"0B25", x"0706", x"037A", x"00BC", x"FEA0", x"FCEE",
		x"FB27", x"F913", x"F69D", x"F3CD", x"F0D8", x"EE33", x"EC34", x"EB30",
		x"EAC9", x"EAA5", x"EADF", x"EC95", x"F0C1", x"F7A3", x"FFDC", x"07D9",
		x"0E38", x"1272", x"149D", x"1501", x"13E3", x"112A", x"0C60", x"058B",
		x"FD5E", x"F56C", x"EF69", x"ED3D", x"EF71", x"F58E", x"FDE7", x"063E",
		x"0CCF", x"1127", x"13B9", x"14D6", x"146F", x"11BF", x"0CB4", x"0587",
		x"FD48", x"F565", x"EF15", x"EB69", x"EA0F", x"EA4A", x"EB00", x"EBF9",
		x"ED89", x"EFD9", x"F26C", x"F48C", x"F55C", x"F475", x"F229", x"EF60",
		x"ECEC", x"EB48", x"EA5D", x"EA10", x"EA86", x"EC44", x"EF97", x"F4B2",
		x"FB9B", x"0374", x"0AF6", x"10B3", x"13D9", x"14BB", x"142C", x"12E1",
		x"1197", x"107D", x"0F6B", x"0E2E", x"0C81", x"0A41", x"0787", x"046C",
		x"00D2", x"FD26", x"FA09", x"F7B3", x"F631", x"F5A9", x"F658", x"F83C",
		x"FB3B", x"FEF4", x"02A5", x"05E1", x"0824", x"0927", x"0876", x"063B",
		x"02BF", x"FEED", x"FB78", x"F8E1", x"F764", x"F701", x"F84A", x"FB7E",
		x"0076", x"06B5", x"0CF4", x"11AB", x"1361", x"115B", x"0BF3", x"043C",
		x"FBE1", x"F45A", x"EEE3", x"EC16", x"EBFD", x"ED92", x"EFD7", x"F1D8",
		x"F2D6", x"F26D", x"F0EE", x"EEDF", x"ECE6", x"EB7E", x"EAE7", x"EB04",
		x"EBBF", x"ECAE", x"ED92", x"EE8C", x"EFC1", x"F18C", x"F3BF", x"F66F",
		x"F98A", x"FD57", x"0161", x"0571", x"08E1", x"0B3D", x"0C13", x"0B1A",
		x"07F0", x"0280", x"FB89", x"F473", x"EF38", x"ECF1", x"ED81", x"EF8A",
		x"F1A9", x"F284", x"F1B8", x"EFC5", x"ED6F", x"EBA6", x"EAB0", x"EA46",
		x"EA58", x"EB6B", x"EE93", x"F458", x"FC42", x"04C0", x"0C24", x"116C",
		x"143A", x"14A5", x"129D", x"0E35", x"07C1", x"FFF4", x"F7EC", x"F120",
		x"ECBD", x"EB6A", x"EC74", x"EE99", x"F10A", x"F319", x"F487", x"F562",
		x"F5C4", x"F5B3", x"F568", x"F496", x"F371", x"F1B8", x"EFB8", x"EDBC",
		x"EC16", x"EB20", x"EAE2", x"EB0E", x"EB85", x"EC0D", x"ECB0", x"ED7A",
		x"EE93", x"F02D", x"F28C", x"F5B1", x"F95D", x"FD57", x"0137", x"04A8",
		x"06F4", x"0781", x"05A2", x"0146", x"FB16", x"F463", x"EF21", x"ECE5",
		x"EDF3", x"F11E", x"F485", x"F6BB", x"F700", x"F566", x"F29D", x"EFAA",
		x"ED59", x"EC0A", x"EB9B", x"EC26", x"EE13", x"F1DC", x"F7A6", x"FEE7",
		x"06BD", x"0DD4", x"1260", x"1344", x"10B3", x"0B42", x"0444", x"FCC4",
		x"F5BE", x"F034", x"ECC8", x"EB8B", x"EBF6", x"EDA5", x"EFE8", x"F265",
		x"F4A1", x"F63E", x"F739", x"F781", x"F75C", x"F68E", x"F581", x"F401",
		x"F222", x"F021", x"EE33", x"ECA1", x"EBB1", x"EB2B", x"EAFE", x"EAE8",
		x"EADD", x"EB08", x"EBB0", x"ED3F", x"F043", x"F54E", x"FC65", x"04B7",
		x"0C6F", x"11C4", x"13F7", x"13C4", x"12BC", x"1257", x"12CF", x"1342",
		x"125E", x"0ECD", x"084E", x"002C", x"F888", x"F346", x"F125", x"F1EB",
		x"F4BA", x"F898", x"FCC7", x"0083", x"0315", x"03A4", x"01A0", x"FD74",
		x"F7F8", x"F27C", x"EE60", x"ECD6", x"EED7", x"F42C", x"FBE5", x"0460",
		x"0BCD", x"1109", x"136B", x"12E4", x"0FF3", x"0BFF", x"089B", x"06EF",
		x"0727", x"08DC", x"0B86", x"0EAD", x"1167", x"132B", x"1404", x"13FC",
		x"1378", x"124E", x"1075", x"0E05", x"0B72", x"090A", x"0718", x"0623",
		x"061F", x"0707", x"08A5", x"0A89", x"0CC1", x"0F1B", x"1178", x"1348",
		x"13A7", x"11CC", x"0D43", x"0688", x"FE9D", x"F71D", x"F12B", x"EDB1",
		x"EC6E", x"ECAA", x"EDD8", x"EFA8", x"F202", x"F4C9", x"F7A4", x"F9CB",
		x"FAC5", x"FA59", x"F888", x"F5F9", x"F320", x"F08E", x"EEA9", x"ED74",
		x"ED0D", x"ECDC", x"ECD1", x"ED25", x"EDFE", x"EF94", x"F214", x"F5B8",
		x"FAB0", x"00E5", x"07B0", x"0DBF", x"11E8", x"1358", x"120A", x"0E9A",
		x"0A48", x"06AE", x"04AC", x"048F", x"05E4", x"085D", x"0B7E", x"0EBC",
		x"119F", x"1389", x"1487", x"14E3", x"14D3", x"1482", x"142E", x"1377",
		x"12B2", x"120B", x"11A3", x"1175", x"11B4", x"125E", x"1348", x"1438",
		x"1482", x"139F", x"1110", x"0C94", x"0636", x"FEA5", x"F730", x"F11B",
		x"ED4F", x"EBAC", x"EB8A", x"EC0F", x"EC6E", x"EC63", x"EBD7", x"EB53",
		x"EB61", x"EC6B", x"EF18", x"F3D1", x"FA6E", x"0219", x"097A", x"0F71",
		x"1319", x"146A", x"13F4", x"128C", x"1151", x"10E5", x"1176", x"12DA",
		x"1464", x"14E4", x"137F", x"10B5", x"0E4A", x"0E0F", x"1011", x"1298",
		x"1347", x"1138", x"0D06", x"085D", x"049C", x"02A0", x"0275", x"03B9",
		x"064A", x"09D2", x"0D9B", x"111C", x"138E", x"1454", x"12B1", x"0E9C",
		x"0826", x"007F", x"F90A", x"F2C4", x"EE73", x"EBF6", x"EAFA", x"EADA",
		x"EB28", x"EB70", x"EBC8", x"EC68", x"EDE7", x"F104", x"F66B", x"FD93",
		x"0565", x"0C59", x"113A", x"13B3", x"13C8", x"1219", x"0F5C", x"0CB0",
		x"0AAD", x"093B", x"07C0", x"0574", x"0212", x"FDCD", x"F8D8", x"F3B8",
		x"EF58", x"ECA3", x"EC98", x"EF87", x"F4FF", x"FC25", x"03DC", x"0B20",
		x"10AD", x"13C8", x"13FB", x"116B", x"0C77", x"05DA", x"FE74", x"F752",
		x"F14D", x"ED5D", x"EBEF", x"ED6F", x"F1AD", x"F7F7", x"FF3D", x"068C",
		x"0CCB", x"116B", x"13C7", x"1370", x"1031", x"0A87", x"0372", x"FBD6",
		x"F4C2", x"EF42", x"EC18", x"EB8D", x"ED9C", x"F251", x"F906", x"011F",
		x"0924", x"0F58", x"12B6", x"1290", x"0F91", x"0AE2", x"069B", x"048F",
		x"055B", x"08D5", x"0D6E", x"1180", x"132F", x"1180", x"0C4D", x"04AD",
		x"FC35", x"F4B3", x"EF4A", x"EC7E", x"EC54", x"EEB1", x"F33C", x"F99C",
		x"00F5", x"0836", x"0E54", x"1256", x"13E8", x"12B2", x"0EF6", x"08EE",
		x"0177", x"F9E1", x"F34D", x"EEA6", x"EC21", x"EC36", x"EEF0", x"F43D",
		x"FB72", x"03A6", x"0B5A", x"10D5", x"12D3", x"1116", x"0CBF", x"07DC",
		x"0488", x"042D", x"0710", x"0C11", x"10ED", x"1329", x"11E8", x"0DC8",
		x"090B", x"05EE", x"05BD", x"0874", x"0CDB", x"10D7", x"126D", x"1075",
		x"0B06", x"0335", x"FAD0", x"F363", x"EE1B", x"EB6E", x"EB8A", x"EE05",
		x"F2D9", x"F99F", x"0190", x"0935", x"0F61", x"12DE", x"136D", x"1144",
		x"0CEB", x"0773", x"01FD", x"FD3B", x"F935", x"F60F", x"F373", x"F17E",
		x"EFEC", x"EE85", x"ED50", x"EC5F", x"EBCF", x"EB82", x"EB19", x"EAD0",
		x"EAEB", x"EBD4", x"EDD8", x"F0CF", x"F525", x"FAD7", x"019B", x"0889",
		x"0E9D", x"1265", x"1337", x"10D6", x"0BC5", x"0527", x"FDDC", x"F6E7",
		x"F120", x"ED45", x"EBCE", x"ED42", x"F1D9", x"F94C", x"0269", x"0B20",
		x"112C", x"13EE", x"142B", x"13C6", x"13BE", x"13FA", x"133F", x"104C",
		x"0AAF", x"0328", x"FB02", x"F478", x"F13D", x"F26E", x"F7CA", x"FFC9",
		x"080D", x"0E8A", x"125B", x"13DC", x"1452", x"1464", x"13FB", x"12A6",
		x"0F57", x"0981", x"01B3", x"F9BE", x"F3BF", x"F14D", x"F2FC", x"F82F",
		x"FF73", x"0750", x"0E1B", x"127D", x"13D1", x"124E", x"0EF3", x"0B36",
		x"0800", x"05BC", x"0416", x"02A8", x"0108", x"FF0B", x"FCC1", x"FA34",
		x"F77A", x"F4C2", x"F24E", x"F05E", x"EED4", x"ED8F", x"EC58", x"EB33",
		x"EA79", x"EA51", x"EABC", x"EB91", x"ECC6", x"EE1E", x"EF88", x"F13B",
		x"F2D8", x"F45A", x"F59A", x"F6E2", x"F8ED", x"FC73", x"0185", x"077C",
		x"0D27", x"113F", x"1258", x"1015", x"0B38", x"05B5", x"01C3", x"0106",
		x"03E0", x"0933", x"0EED", x"12A6", x"12DD", x"102E", x"0C28", x"0922",
		x"08A0", x"0AC1", x"0EA8", x"11D9", x"1278", x"0F4B", x"08E2", x"009A",
		x"F853", x"F1A5", x"ED55", x"EB83", x"EC45", x"EF72", x"F4ED", x"FC20",
		x"03ED", x"0B23", x"105A", x"12A3", x"11A2", x"0DE8", x"08E5", x"040E",
		x"0067", x"FE9B", x"FE9A", x"003A", x"0300", x"062C", x"0957", x"0C0C",
		x"0E0F", x"0F25", x"0F60", x"0EC4", x"0D49", x"0ADC", x"0782", x"031E",
		x"FE2D", x"F915", x"F42D", x"EFFE", x"ED15", x"EC45", x"EE73", x"F365",
		x"FA72", x"0278", x"0A26", x"100A", x"1338", x"1348", x"10A2", x"0C3C",
		x"0686", x"0081", x"FAF4", x"F64F", x"F2A9", x"EFF5", x"EE15", x"ECDB",
		x"EC38", x"EBFF", x"EC18", x"ECE1", x"EE6A", x"F0E5", x"F3FA", x"F719",
		x"F99B", x"FA8B", x"F929", x"F5B8", x"F165", x"EE35", x"EDB7", x"F0C6",
		x"F671", x"FC9C", x"00AF", x"00FD", x"FD46", x"F719", x"F12B", x"EDD4",
		x"EE19", x"F11B", x"F48B", x"F640", x"F538", x"F1E4", x"EE72", x"ED85",
		x"F016", x"F5ED", x"FCAF", x"022C", x"04E9", x"04C9", x"025D", x"FE91",
		x"FA6B", x"F68B", x"F3D0", x"F251", x"F241", x"F34E", x"F574", x"F89D",
		x"FC59", x"FFE0", x"02B5", x"045C", x"04AA", x"0389", x"0142", x"FE1F",
		x"FADE", x"F7E7", x"F55D", x"F38E", x"F28F", x"F298", x"F385", x"F539",
		x"F768", x"FA23", x"FD58", x"00E4", x"0480", x"07BC", x"0AC5", x"0DA4",
		x"102F", x"1220", x"1356", x"13C0", x"1413", x"1427", x"13FA", x"135A",
		x"1210", x"1033", x"0DEE", x"0B8D", x"0972", x"0819", x"07E9", x"08D4",
		x"0AB6", x"0D19", x"0F9A", x"11CF", x"137F", x"149F", x"152D", x"1569",
		x"1553", x"150E", x"148C", x"13B5", x"1250", x"0FE8", x"0C15", x"067B",
		x"FF3B", x"F79D", x"F117", x"ED02", x"EBD7", x"ED51", x"F091", x"F475",
		x"F81F", x"FB46", x"FE10", x"007C", x"02D1", x"04CA", x"0667", x"0803",
		x"0990", x"0B36", x"0CD8", x"0E81", x"1049", x"1226", x"13CD", x"147D",
		x"13E5", x"1167", x"0CD5", x"068E", x"FF4C", x"F805", x"F1C2", x"EDC4",
		x"ED82", x"F144", x"F85B", x"00CC", x"0887", x"0E35", x"11AC", x"135C",
		x"137C", x"11D0", x"0E5D", x"08D8", x"0199", x"F984", x"F239", x"EDAD",
		x"ED35", x"F134", x"F8B5", x"01CA", x"0A25", x"1045", x"13D5", x"1568",
		x"15B1", x"149E", x"11B1", x"0C99", x"0580", x"FD71", x"F5A3", x"EF6F",
		x"EBBD", x"EB30", x"ED9E", x"F2B6", x"F9C7", x"01DB", x"09A6", x"0FEE",
		x"13DB", x"157F", x"1577", x"14FB", x"14C0", x"14CD", x"1471", x"12EC",
		x"0FC8", x"0B36", x"0571", x"FEC5", x"F7EC", x"F1FF", x"EDDE", x"EC7A",
		x"EDAF", x"F0C9", x"F4E0", x"F8BB", x"FBFA", x"FE8F", x"00BD", x"02E4",
		x"04D9", x"06BE", x"08A1", x"0A94", x"0CA2", x"0E9D", x"106D", x"11EF",
		x"130E", x"13EA", x"149F", x"1505", x"14C8", x"13AB", x"11EE", x"0FF7",
		x"0E75", x"0DB0", x"0DEE", x"0F5C", x"1185", x"1371", x"13D0", x"1167",
		x"0BFF", x"0440", x"FBB9", x"F416", x"EECD", x"EC6B", x"ECBF", x"EF58",
		x"F3A0", x"F989", x"00B2", x"0868", x"0EEA", x"1276", x"11FF", x"0DD8",
		x"07A0", x"0116", x"FBE7", x"F909", x"F967", x"FCDC", x"029D", x"0937",
		x"0F04", x"1291", x"1316", x"10B9", x"0C37", x"06BB", x"0141", x"FC74",
		x"F8A7", x"F640", x"F574", x"F680", x"F952", x"FE17", x"0459", x"0B30",
		x"10C5", x"137B", x"134C", x"111C", x"0EF9", x"0E4E", x"0F9D", x"11D8",
		x"1313", x"1193", x"0C8F", x"0518", x"FD0C", x"F671", x"F202", x"EFAA",
		x"EEAC", x"EE72", x"EE38", x"ED67", x"EC45", x"EBA0", x"ECDA", x"F0D5",
		x"F765", x"FF44", x"0704", x"0D6D", x"11DE", x"1477", x"156D", x"157F",
		x"1520", x"14B7", x"13FE", x"12A1", x"107B", x"0D7C", x"09E8", x"05F0",
		x"01D1", x"FDD4", x"FA5D", x"F774", x"F5B1", x"F597", x"F7AC", x"FC23",
		x"0283", x"0993", x"0F98", x"12FF", x"135C", x"11A2", x"0F99", x"0EEF",
		x"1022", x"1224", x"1317", x"112A", x"0BC0", x"03FE", x"FBF2", x"F576",
		x"F15A", x"EF47", x"EE64", x"EDE4", x"ED47", x"EC8B", x"EB8D", x"EB4C",
		x"ECAC", x"F080", x"F6F3", x"FEEC", x"06F1", x"0DB4", x"1248", x"14A5",
		x"1569", x"152E", x"1481", x"1376", x"11F0", x"0FA1", x"0D5F", x"0B97",
		x"0B00", x"0BBC", x"0D77", x"0FDB", x"122E", x"1405", x"1505", x"1582",
		x"153F", x"1387", x"0F83", x"08E5", x"00B6", x"F899", x"F1DC", x"ED4D",
		x"EAF2", x"EAB2", x"EC2B", x"EFA2", x"F535", x"FCF2", x"056B", x"0D18",
		x"1257", x"14C0", x"14F8", x"13F8", x"12C7", x"11AF", x"10A8", x"0F88",
		x"0E1F", x"0C28", x"09C0", x"06F6", x"03F7", x"00BE", x"FD8A", x"FAAE",
		x"F888", x"F799", x"F7F0", x"F98D", x"FC02", x"FF58", x"02E1", x"0648",
		x"0919", x"0AD4", x"0B31", x"09EE", x"0735", x"036E", x"FF10", x"FB0A",
		x"F803", x"F6F1", x"F851", x"FC7A", x"0304", x"0A4F", x"103C", x"1302",
		x"124C", x"0FBF", x"0DB3", x"0D6F", x"0F4A", x"11C5", x"12F2", x"1142",
		x"0C71", x"057F", x"FE94", x"F979", x"F715", x"F749", x"F976", x"FCD1",
		x"00CC", x"04DA", x"08AF", x"0C0F", x"0E9B", x"107D", x"11D5", x"12CD",
		x"13AD", x"147F", x"14FE", x"1521", x"14D4", x"1427", x"12DF", x"10EC",
		x"0EAB", x"0C6B", x"0ADA", x"0A02", x"0A02", x"0AD0", x"0C61", x"0E72",
		x"10A7", x"127A", x"13BB", x"1477", x"1497", x"1459", x"1386", x"11FE",
		x"0FAB", x"0CB1", x"0A00", x"088A", x"0917", x"0BC1", x"0F46", x"1222",
		x"129C", x"0FE4", x"0A6B", x"03F8", x"FED1", x"FC92", x"FE33", x"031E",
		x"099B", x"0F6C", x"1288", x"123D", x"0EFF", x"09EB", x"046D", x"FFAB",
		x"FC80", x"FA7F", x"F908", x"F7A3", x"F5ED", x"F412", x"F240", x"F075",
		x"EED0", x"ED57", x"EC26", x"EB65", x"EB01", x"EB13", x"EB7F", x"EC64",
		x"EDA8", x"EF6B", x"F180", x"F3AE", x"F5AA", x"F70F", x"F794", x"F6ED",
		x"F52A", x"F29B", x"EFCA", x"ED8B", x"EBE9", x"EB10", x"EB10", x"ECA1",
		x"F095", x"F742", x"FF9C", x"0803", x"0EC7", x"1355", x"15BC", x"1642",
		x"14E5", x"1151", x"0BA5", x"041C", x"FBE7", x"F464", x"EED7", x"EC16",
		x"EC64", x"EF5A", x"F48C", x"FB7C", x"038F", x"0B58", x"1141", x"1439",
		x"1443", x"1277", x"1042", x"0E9E", x"0D8E", x"0CC6", x"0BA0", x"09CD",
		x"0740", x"041B", x"0079", x"FC7F", x"F8BB", x"F5B8", x"F3AA", x"F2C7",
		x"F2C4", x"F3AD", x"F549", x"F796", x"FA51", x"FD11", x"FF93", x"01A3",
		x"032C", x"041C", x"0445", x"03BB", x"027E", x"0076", x"FD9D", x"F9A9",
		x"F4E5", x"F060", x"ED5C", x"ED3C", x"F005", x"F57B", x"FC55", x"0351",
		x"08C6", x"0B3D", x"0A2C", x"05A0", x"FEDE", x"F793", x"F15A", x"ED8D",
		x"ECA6", x"EE01", x"F02D", x"F1A1", x"F13D", x"EF6B", x"ED4D", x"EBC3",
		x"EB44", x"EB6E", x"EC09", x"ECE2", x"EDC3", x"EEB4", x"EF8E", x"F0CA",
		x"F2C6", x"F634", x"FB3D", x"01C0", x"08C9", x"0EE2", x"12CA", x"13B4",
		x"11B2", x"0E18", x"0A4E", x"0788", x"066A", x"0769", x"09E7", x"0D1E",
		x"1050", x"12A1", x"13EF", x"1451", x"13C6", x"123B", x"0F9A", x"0C14",
		x"084C", x"0547", x"0416", x"0575", x"0938", x"0DFA", x"11BF", x"1291",
		x"0FD6", x"0A78", x"049E", x"00AC", x"002F", x"038F", x"0943", x"0EEE",
		x"123E", x"1248", x"0F34", x"0AB1", x"067B", x"0412", x"03EE", x"05CC",
		x"08DA", x"0C34", x"0F75", x"121C", x"13F6", x"14EF", x"1515", x"14BF",
		x"140B", x"133F", x"1276", x"11CF", x"1153", x"114F", x"11D5", x"12B2",
		x"13B4", x"148C", x"1534", x"1537", x"14CA", x"144F", x"142C", x"1467",
		x"14AB", x"1496", x"13E7", x"12B1", x"117D", x"110D", x"1199", x"12E2",
		x"140E", x"148F", x"1456", x"13FA", x"13E4", x"1440", x"1490", x"13F9",
		x"1171", x"0C83", x"0570", x"FD63", x"F5F4", x"F07B", x"ED68", x"EC74",
		x"ECCB", x"EDEB", x"EFE5", x"F294", x"F5F3", x"F970", x"FD05", x"0021",
		x"02E8", x"0564", x"07C2", x"0A05", x"0C44", x"0E57", x"1020", x"11CB",
		x"1310", x"13FC", x"148A", x"14EE", x"1502", x"14BF", x"1418", x"1309",
		x"118D", x"0FCC", x"0DA0", x"0B34", x"08C6", x"06DE", x"05A0", x"04F9",
		x"04D3", x"0530", x"0623", x"079B", x"0975", x"0BCD", x"0EAE", x"11B6",
		x"13B1", x"1322", x"0F68", x"0909", x"016F", x"F9D5", x"F3BD", x"F005",
		x"EEF9", x"F062", x"F429", x"F9F6", x"015A", x"0958", x"0FDE", x"1341",
		x"1274", x"0DE4", x"06DE", x"FEE6", x"F766", x"F147", x"ED31", x"EB85",
		x"EBF0", x"EDA2", x"EFD8", x"F1CA", x"F357", x"F4C6", x"F658", x"F883",
		x"FBBB", x"0045", x"0609", x"0C30", x"10E3", x"12E4", x"1155", x"0D35",
		x"0836", x"0461", x"02CE", x"03A4", x"0661", x"09F0", x"0D7E", x"100D",
		x"1185", x"11B4", x"106A", x"0D64", x"089B", x"0212", x"FA91", x"F376",
		x"EE50", x"ECC0", x"EF3E", x"F57E", x"FE08", x"06E1", x"0DFE", x"1277",
		x"1477", x"14E4", x"14F2", x"1503", x"1496", x"128E", x"0E58", x"0798",
		x"FF67", x"F753", x"F0DD", x"ECC4", x"EAE9", x"EA6F", x"EAAA", x"EB2A",
		x"EBC1", x"EC6B", x"ED44", x"EE47", x"EF66", x"F0CC", x"F205", x"F387",
		x"F55F", x"F7FF", x"FBEA", x"00FC", x"06E2", x"0CA1", x"10F0", x"12F8",
		x"1231", x"0ED7", x"0A08", x"0540", x"01AF", x"0032", x"006A", x"0217",
		x"04BE", x"081A", x"0BD1", x"0F79", x"1266", x"1355", x"118C", x"0CA2",
		x"0587", x"FD91", x"F650", x"F13A", x"EF42", x"F114", x"F669", x"FE3A",
		x"068B", x"0DA5", x"1276", x"14FD", x"15BE", x"15B1", x"14FB", x"136A",
		x"0FDC", x"09FF", x"0215", x"F9F8", x"F341", x"EEEE", x"ECF9", x"ECCD",
		x"ED81", x"EF30", x"F1DE", x"F5C8", x"FAB4", x"005F", x"0652", x"0BF9",
		x"10A3", x"1365", x"1388", x"10DD", x"0C0B", x"05FD", x"FFE8", x"FA73",
		x"F61C", x"F33D", x"F170", x"F065", x"EFC8", x"EF8A", x"EFD1", x"F063",
		x"F144", x"F25D", x"F3EB", x"F605", x"F8E4", x"FC65", x"007E", x"04A9",
		x"0899", x"0BED", x"0E9E", x"109A", x"11DF", x"1262", x"11CB", x"0FE5",
		x"0C8F", x"07AC", x"013E", x"FA09", x"F32F", x"EE2E", x"EC72", x"EE9A",
		x"F42E", x"FBC6", x"03BE", x"0AC2", x"100A", x"135D", x"14A0", x"13F9",
		x"11C5", x"0E85", x"0ACF", x"06F4", x"03BF", x"01B6", x"01C3", x"03A6",
		x"0757", x"0BED", x"105F", x"1350", x"13AC", x"1131", x"0C79", x"066F",
		x"FFFF", x"F9E4", x"F4AB", x"F0C7", x"EE1B", x"EC99", x"EC01", x"EC47",
		x"EDBF", x"F156", x"F75C", x"FF3F", x"0768", x"0E18", x"1297", x"14F8",
		x"1612", x"1615", x"152C", x"130E", x"0EF6", x"08BD", x"00B2", x"F88D",
		x"F1E9", x"EDD7", x"EC1A", x"EBEA", x"ECBA", x"EE53", x"F0E8", x"F474",
		x"F90C", x"FEA0", x"04C6", x"0AEE", x"1018", x"133E", x"13BB", x"1182",
		x"0D29", x"079F", x"0210", x"FCEC", x"F90A", x"F698", x"F53B", x"F465",
		x"F373", x"F234", x"F077", x"EE90", x"ECF4", x"EBC2", x"EB4B", x"EB10",
		x"EB30", x"EB55", x"EB7C", x"EB84", x"EB4D", x"EB24", x"EB42", x"EBE4",
		x"ECC3", x"ED85", x"EDBE", x"ED13", x"EC14", x"EBBA", x"ED77", x"F1F8",
		x"F911", x"01A2", x"09CF", x"1020", x"13AA", x"142E", x"11DF", x"0D4B",
		x"0723", x"0038", x"F92E", x"F2C1", x"EE59", x"ECDD", x"EEFA", x"F458",
		x"FBAE", x"030F", x"092C", x"0D35", x"0F02", x"0F23", x"0E0B", x"0C5E",
		x"0A21", x"075B", x"03F3", x"0007", x"FC0B", x"F82D", x"F478", x"F11A",
		x"EE6A", x"EC91", x"EB93", x"EB61", x"EC5F", x"EF89", x"F55D", x"FD40",
		x"0583", x"0CC6", x"11D1", x"14B8", x"15BB", x"1598", x"14BB", x"12BE",
		x"0EEB", x"08A8", x"009B", x"F809", x"F12F", x"ECE5", x"EB65", x"EBC9",
		x"ED26", x"EE98", x"EFC3", x"F041", x"EFE3", x"EEA3", x"ED1F", x"EC50",
		x"ED41", x"F0BB", x"F698", x"FE12", x"0592", x"0B6F", x"0ECC", x"0F94",
		x"0E48", x"0B5D", x"077E", x"02F4", x"FEB6", x"FBC9", x"FAFB", x"FC29",
		x"FF59", x"037C", x"07CD", x"0B61", x"0DD0", x"0EAA", x"0D87", x"09EB",
		x"03F2", x"FC4F", x"F4E0", x"EF55", x"EC7A", x"EC47", x"EDBE", x"EF86",
		x"F07C", x"F030", x"EEE5", x"ED28", x"EBC4", x"EB10", x"EB23", x"EBE3",
		x"ED4B", x"EED9", x"F046", x"F199", x"F2D2", x"F460", x"F67B", x"F92C",
		x"FC6B", x"001F", x"03AD", x"06E4", x"0992", x"0BA4", x"0D09", x"0D90",
		x"0D27", x"0BCF", x"09AD", x"06F7", x"0411", x"0136", x"FECB", x"FD2A",
		x"FC22", x"FBC5", x"FC08", x"FD06", x"FEC5", x"0172", x"04FC", x"0973",
		x"0E22", x"11DC", x"1336", x"1191", x"0CF8", x"0669", x"FF66", x"F96D",
		x"F5D9", x"F5AE", x"F8EB", x"FECE", x"061A", x"0CDB", x"117E", x"1321",
		x"11CC", x"0E61", x"0A2B", x"0632", x"030A", x"00D4", x"FF42", x"FDB9",
		x"FC08", x"F9EE", x"F7D3", x"F5DA", x"F414", x"F282", x"F0F5", x"EF46",
		x"ED66", x"EBD7", x"EBA5", x"ED98", x"F1FE", x"F88F", x"0046", x"07EE",
		x"0E89", x"1314", x"1549", x"1585", x"1471", x"1288", x"0FD3", x"0CA5",
		x"09A5", x"0806", x"08B1", x"0B9C", x"0F62", x"11D1", x"1149", x"0D34",
		x"06C6", x"0045", x"FC31", x"FC3D", x"009A", x"0793", x"0E8A", x"129D",
		x"12E1", x"102B", x"0D0B", x"0BA3", x"0CAF", x"0F6C", x"11E8", x"1248",
		x"0F3B", x"0924", x"01E9", x"FBC6", x"F80A", x"F714", x"F87E", x"FB70",
		x"FF46", x"039A", x"07D3", x"0B73", x"0E40", x"1047", x"11B9", x"12D2",
		x"13B6", x"1471", x"1505", x"1569", x"1531", x"147B", x"1328", x"1127",
		x"0ED5", x"0CA9", x"0AFA", x"0A23", x"0A0C", x"0A74", x"0B3A", x"0C68",
		x"0E24", x"100D", x"120A", x"13B0", x"14EB", x"1564", x"14EF", x"13A0",
		x"11BB", x"0F9E", x"0DDC", x"0CF3", x"0D65", x"0F22", x"116C", x"12E7",
		x"123F", x"0E96", x"086E", x"0129", x"FAE5", x"F798", x"F80C", x"FC25",
		x"02A7", x"09A2", x"0F3D", x"1202", x"11A6", x"0EBF", x"0ABF", x"06CF",
		x"03CE", x"01FD", x"00D4", x"FFCB", x"FDC6", x"FA64", x"F5D2", x"F110",
		x"ED73", x"EC54", x"EE25", x"F2A3", x"F8EC", x"FF89", x"0585", x"0A85",
		x"0E66", x"1155", x"133F", x"143D", x"14CF", x"151C", x"152F", x"1500",
		x"145E", x"1309", x"10D9", x"0E3B", x"0B8E", x"0A14", x"0A41", x"0C4D",
		x"0F57", x"11F4", x"12A6", x"1058", x"0B2B", x"048C", x"FE88", x"FB07",
		x"FAE1", x"FE16", x"03A7", x"0A3B", x"0FDF", x"12CC", x"11EB", x"0CF4",
		x"053C", x"FC96", x"F4F3", x"EF82", x"EC82", x"EC09", x"ED9B", x"F0D5",
		x"F52B", x"F9F6", x"FE67", x"022A", x"0541", x"07AB", x"094F", x"0A0D",
		x"09D7", x"087A", x"0682", x"03BB", x"0065", x"FCDF", x"F9CF", x"F7A5",
		x"F6BE", x"F743", x"F91A", x"FC02", x"FF69", x"0304", x"0640", x"0884",
		x"0951", x"07F9", x"0454", x"FEE5", x"F8A4", x"F284", x"EE28", x"ECB7",
		x"EEE9", x"F499", x"FCB0", x"054E", x"0CC2", x"11E9", x"143F", x"13EF",
		x"11BF", x"0EF4", x"0D00", x"0C77", x"0D58", x"0F19", x"112E", x"1314",
		x"1472", x"1519", x"1569", x"1574", x"1542", x"14B1", x"13AE", x"121B",
		x"100C", x"0D94", x"0AAE", x"076F", x"03B3", x"FF98", x"FB92", x"F826",
		x"F5F8", x"F528", x"F62A", x"F94C", x"FEA2", x"0582", x"0C63", x"1163",
		x"1373", x"12AB", x"102F", x"0DA8", x"0C65", x"0CD4", x"0EB6", x"1127",
		x"1341", x"14BA", x"155D", x"1575", x"152D", x"1493", x"1387", x"11CF",
		x"0FC0", x"0DFB", x"0D13", x"0D8F", x"0F31", x"1162", x"131C", x"1309",
		x"1048", x"0AC1", x"0373", x"FBDF", x"F54B", x"F070", x"ED77", x"EBF8",
		x"EB3A", x"EAD2", x"EA9C", x"EA7C", x"EA8F", x"EA97", x"EA98", x"EACE",
		x"EB86", x"ECAB", x"EE2B", x"EFF3", x"F221", x"F4E2", x"F843", x"FBE9",
		x"FF9F", x"02F1", x"058B", x"0732", x"07E4", x"0796", x"0605", x"033C",
		x"FF7C", x"FBA0", x"F854", x"F630", x"F55D", x"F624", x"F915", x"FE38",
		x"04C4", x"0B62", x"10BC", x"1361", x"1302", x"0FEE", x"0B1B", x"05D2",
		x"011F", x"FD3E", x"FA57", x"F8AB", x"F80A", x"F8E6", x"FB5C", x"FFA8",
		x"0541", x"0B58", x"1058", x"12FC", x"1293", x"0F4C", x"0A37", x"04E0",
		x"0076", x"FD56", x"FB3B", x"F9CA", x"F884", x"F6EC", x"F508", x"F2B0",
		x"F04D", x"EE1F", x"EC7A", x"EB56", x"EAA7", x"EA23", x"E9ED", x"EA48",
		x"EBD3", x"EF2C", x"F48F", x"FBCC", x"03C7", x"0B5B", x"1115", x"1470",
		x"158C", x"153B", x"148C", x"13C1", x"12FF", x"11FD", x"105B", x"0DAA",
		x"0982", x"03E9", x"FD50", x"F6B4", x"F11E", x"ED5C", x"EC5E", x"EEA6",
		x"F42F", x"FC20", x"04D3", x"0CB3", x"1243", x"14CB", x"14B4", x"12DE",
		x"10EB", x"0FD8", x"1029", x"1182", x"132D", x"1482", x"1538", x"158C",
		x"15A3", x"157A", x"148E", x"1220", x"0D99", x"0690", x"FE14", x"F59B",
		x"EF17", x"EC2F", x"ECCA", x"F04F", x"F590", x"FBE9", x"02BC", x"099D",
		x"0F93", x"1351", x"13C4", x"1073", x"0A01", x"01F1", x"FA10", x"F3B0",
		x"EF36", x"EC9A", x"EB7D", x"EB74", x"EC5A", x"EDDE", x"EFC7", x"F1FF",
		x"F42C", x"F63A", x"F7A1", x"F839", x"F7E0", x"F6C4", x"F511", x"F2DB",
		x"F033", x"ED8D", x"EBF9", x"EC63", x"EFA4", x"F5A8", x"FD4F", x"0540",
		x"0BFF", x"10BB", x"1344", x"1370", x"1152", x"0CCE", x"0647", x"FE3E",
		x"F638", x"EFE4", x"EC4F", x"EBD9", x"ED9A", x"F058", x"F2E3", x"F52B",
		x"F707", x"F867", x"F921", x"F8D8", x"F771", x"F541", x"F292", x"F019",
		x"EE49", x"ED14", x"EC3C", x"EC15", x"ED46", x"F0B2", x"F6B9", x"FE89",
		x"06BD", x"0E08", x"1305", x"158A", x"15FB", x"1571", x"1502", x"14A4",
		x"13F4", x"12B9", x"113B", x"1040", x"1097", x"11F3", x"1332", x"129F",
		x"0F63", x"0924", x"0180", x"FA1D", x"F494", x"F1AE", x"F146", x"F2C1",
		x"F57C", x"F92C", x"FD03", x"00A0", x"034A", x"0457", x"039D", x"0158",
		x"FE22", x"FAAC", x"F749", x"F46C", x"F274", x"F185", x"F19A", x"F2A9",
		x"F486", x"F6E3", x"F9C0", x"FCDB", x"0024", x"0359", x"064F", x"08D5",
		x"0B16", x"0D05", x"0ED7", x"1071", x"11E9", x"1332", x"141A", x"14B2",
		x"14FF", x"1516", x"14CE", x"1453", x"1366", x"121E", x"107C", x"0E7A",
		x"0BE5", x"08E1", x"05D7", x"0308", x"00E1", x"FF3C", x"FE2D", x"FDA3",
		x"FDF4", x"FF30", x"011D", x"03B1", x"0695", x"09FC", x"0DB3", x"1123",
		x"1366", x"13D3", x"1223", x"0E07", x"07C4", x"0028", x"F86A", x"F1D5",
		x"ED81", x"EC02", x"ED64", x"F15F", x"F737", x"FE25", x"0557", x"0BE4",
		x"10F4", x"1388", x"12FA", x"0F54", x"0963", x"0252", x"FB22", x"F4D4",
		x"F03C", x"ED67", x"EC06", x"EB73", x"EB30", x"EAE9", x"EA9F", x"EAC5",
		x"EC3E", x"F018", x"F69E", x"FF2E", x"07FC", x"0EE2", x"1318", x"1526",
		x"15E1", x"15AF", x"145C", x"1129", x"0BDF", x"04DB", x"FCE7", x"F598",
		x"F060", x"EE33", x"EF0A", x"F271", x"F7F9", x"FF36", x"073C", x"0E52",
		x"125A", x"1230", x"0D97", x"05BF", x"FCC5", x"F4BD", x"EF16", x"EBFA",
		x"EABE", x"EA72", x"EA81", x"EB01", x"EC8F", x"F031", x"F653", x"FE8A",
		x"0724", x"0E58", x"12D8", x"14D5", x"151D", x"1498", x"13F7", x"136C",
		x"1316", x"12D7", x"12AF", x"1298", x"12B8", x"1306", x"137D", x"1409",
		x"1456", x"1421", x"12EE", x"1003", x"0B1F", x"0450", x"FCAA", x"F563",
		x"EFE2", x"EC9C", x"EBBC", x"ECC3", x"EED6", x"F10C", x"F2D0", x"F425",
		x"F55F", x"F722", x"FA0E", x"FE40", x"03E7", x"0A3E", x"0FC9", x"12D4",
		x"1254", x"0EC9", x"09C6", x"055F", x"0301", x"0348", x"05D4", x"0989",
		x"0D59", x"106F", x"1270", x"131E", x"119C", x"0D8F", x"06EE", x"FEC6",
		x"F6D8", x"F0C4", x"ED27", x"EB78", x"EB0A", x"EAE8", x"EB19", x"EC79",
		x"EFE6", x"F606", x"FE38", x"06D6", x"0E00", x"125C", x"1353", x"10E4",
		x"0BA0", x"048E", x"FD25", x"F6AE", x"F1DD", x"EE77", x"EC36", x"EAF6",
		x"EA97", x"EAE4", x"EB61", x"EC15", x"ECE4", x"EE06", x"EF5B", x"F0DA",
		x"F289", x"F44B", x"F663", x"F88F", x"FB20", x"FDDC", x"0140", x"050D",
		x"08FC", x"0CA3", x"0F6E", x"1122", x"11D9", x"119B", x"1047", x"0D1D",
		x"082B", x"01AF", x"FA86", x"F3D2", x"EED1", x"ECA5", x"EE39", x"F381",
		x"FB93", x"04B5", x"0CAB", x"11D7", x"1446", x"14D6", x"14A7", x"1481",
		x"13FA", x"1219", x"0DE8", x"073F", x"FF22", x"F793", x"F229", x"F006",
		x"F153", x"F5BA", x"FC78", x"0446", x"0B9F", x"1121", x"137C", x"12A0",
		x"0F4D", x"0AEF", x"06B6", x"0356", x"0102", x"FFB4", x"FFA9", x"0143",
		x"049F", x"093E", x"0E3F", x"11D7", x"12ED", x"10F9", x"0CF1", x"0805",
		x"03DD", x"0180", x"017D", x"037E", x"06C9", x"0A79", x"0DD7", x"109B",
		x"129D", x"13CD", x"1474", x"14DD", x"14F1", x"14E5", x"1493", x"13C7",
		x"11CA", x"0DDC", x"07CD", x"001C", x"F811", x"F177", x"ED51", x"EBA6",
		x"EBA2", x"EC79", x"ED4A", x"ED5F", x"ECC6", x"EBBE", x"EAEE", x"EAE9",
		x"EBDB", x"ED5E", x"EED7", x"F006", x"F0B0", x"F129", x"F1E3", x"F393",
		x"F6BB", x"FB78", x"01B8", x"08E0", x"0F33", x"12D9", x"12D4", x"0F6D",
		x"0AB3", x"073E", x"06D3", x"0947", x"0D6C", x"114E", x"12F7", x"1198",
		x"0D66", x"07AF", x"024B", x"FE9A", x"FCFA", x"FD52", x"FF3F", x"023A",
		x"062D", x"0AE7", x"0F88", x"12E3", x"13BF", x"117B", x"0C59", x"0575",
		x"FE0E", x"F784", x"F2F2", x"F194", x"F3CD", x"F95C", x"00E9", x"08A2",
		x"0ED2", x"129D", x"13B5", x"12C8", x"1170", x"10D2", x"1183", x"12D9",
		x"13DF", x"1439", x"1428", x"1402", x"141D", x"146A", x"149E", x"1487",
		x"1409", x"1304", x"11FB", x"116D", x"11EE", x"1315", x"13BA", x"1236",
		x"0DED", x"0708", x"FF2C", x"F7B0", x"F1D2", x"EDF5", x"EBC9", x"EAF2",
		x"EAD5", x"EB1B", x"EB6A", x"EB85", x"EB83", x"EB4E", x"EB04", x"EABB",
		x"EACD", x"EB62", x"EC73", x"ED84", x"EE58", x"EE87", x"EE01", x"ED22",
		x"EC15", x"EB5A", x"EB1F", x"EB44", x"EB6E", x"EB91", x"EB80", x"EB53",
		x"EB50", x"EBCA", x"ECCE", x"EDF6", x"EE9B", x"EE35", x"ED0E", x"EBE8",
		x"EBDD", x"EE06", x"F2CE", x"F9F9", x"021F", x"09AF", x"0F22", x"1277",
		x"1417", x"14E3", x"1528", x"1546", x"1518", x"14E5", x"14D7", x"1502",
		x"1523", x"1525", x"14E9", x"147A", x"138B", x"120F", x"101D", x"0DFF",
		x"0BF7", x"09ED", x"07CB", x"05AF", x"03B0", x"0199", x"FF11", x"FC07",
		x"F891", x"F4F2", x"F197", x"EECD", x"ECC8", x"EBC1", x"EBD9", x"ECEB",
		x"EF2D", x"F2F9", x"F8B2", x"FFD9", x"0782", x"0E4A", x"12BB", x"147B",
		x"1388", x"10E1", x"0D7B", x"0A3C", x"07E2", x"066E", x"0634", x"0749",
		x"0983", x"0C9E", x"0FFC", x"129F", x"1379", x"117E", x"0CA1", x"0535",
		x"FC99", x"F473", x"EE7E", x"EBB8", x"EC0B", x"EF02", x"F3E7", x"F9A9",
		x"FFA6", x"055C", x"0A6D", x"0E62", x"1166", x"1338", x"13FF", x"143B",
		x"140A", x"1304", x"1072", x"0BC3", x"051B", x"FD2F", x"F582", x"EF8A",
		x"EC44", x"EBB4", x"ECE2", x"EE92", x"EFE6", x"F092", x"F0EB", x"F1CC",
		x"F3FF", x"F821", x"FE34", x"0550", x"0C4E", x"118C", x"1397", x"123C",
		x"0EDE", x"0BCB", x"0ADF", x"0CA5", x"0FC9", x"128F", x"12FD", x"1032",
		x"0ABC", x"0416", x"FE0C", x"F9DA", x"F822", x"F8AE", x"FB2C", x"FF00",
		x"03B6", x"08B2", x"0D5D", x"1139", x"13B1", x"146C", x"12DC", x"0EF8",
		x"08F5", x"019C", x"F9C4", x"F29D", x"EDB0", x"EC20", x"EDF2", x"F268",
		x"F858", x"FEBF", x"04EE", x"0A80", x"0F03", x"1225", x"1419", x"14F6",
		x"151D", x"14F8", x"1502", x"151E", x"1535", x"14E0", x"1434", x"1323",
		x"11D4", x"106D", x"0F40", x"0F25", x"1028", x"11EC", x"13AD", x"1429",
		x"1262", x"0DB0", x"067E", x"FDEB", x"F59C", x"EF7E", x"ED10", x"EED4",
		x"F3F2", x"FADA", x"0182", x"06B7", x"096E", x"08E4", x"04F2", x"FE78",
		x"F726", x"F116", x"ED8A", x"ECE0", x"EE50", x"F080", x"F21D", x"F230",
		x"F0BD", x"EE6A", x"EC7B", x"EB44", x"EACB", x"EA95", x"EA85", x"EAC7",
		x"EBB9", x"ED71", x"EF7D", x"F15A", x"F22B", x"F18F", x"EFD2", x"ED88",
		x"EC62", x"ED88", x"F1CC", x"F891", x"0009", x"065D", x"0A5C", x"0BFA",
		x"0BBE", x"0A0D", x"0744", x"03BE", x"FFC5", x"FBE5", x"F841", x"F511",
		x"F239", x"EFCF", x"EE17", x"ED00", x"EC54", x"EBD3", x"EB61", x"EB1F",
		x"EB37", x"EC16", x"EDAF", x"EFBE", x"F20A", x"F3F8", x"F55D", x"F5F3",
		x"F56D", x"F3D6", x"F18B", x"EF18", x"ED1E", x"EBE1", x"EB34", x"EAFA",
		x"EAF7", x"EB1D", x"EB58", x"EBAA", x"EC99", x"EE40", x"F0F8", x"F531",
		x"FAFC", x"01E8", x"0935", x"0F52", x"12EF", x"13B4", x"11FF", x"0F1F",
		x"0C52", x"0AC3", x"0AD9", x"0C5A", x"0E94", x"10FF", x"12EB", x"13F7",
		x"1467", x"1449", x"13FD", x"13B1", x"12EA", x"11A1", x"0FAB", x"0D71",
		x"0B41", x"093B", x"0788", x"0607", x"0498", x"02ED", x"00A8", x"FD6F",
		x"F92E", x"F44C", x"EFC8", x"ECFA", x"ECFB", x"EFC9", x"F4BF", x"FACE",
		x"00E7", x"05C6", x"08E9", x"0A3B", x"0A00", x"08A7", x"064E", x"02B5",
		x"FD9F", x"F798", x"F1E0", x"EDE9", x"ECCF", x"EEF1", x"F3B9", x"F9D0",
		x"FFBA", x"0414", x"05B6", x"046F", x"0095", x"FAF4", x"F4E2", x"EFBE",
		x"ED81", x"EF23", x"F4FB", x"FD4B", x"061C", x"0D5D", x"11FA", x"13BD",
		x"134D", x"1181", x"0F25", x"0CCF", x"0B2F", x"0AA5", x"0B71", x"0D66",
		x"0FFF", x"1299", x"1453", x"1462", x"124D", x"0DCD", x"0792", x"0059",
		x"F91E", x"F2E4", x"EE2E", x"EB90", x"EAFD", x"EC2E", x"EE9D", x"F15A",
		x"F39B", x"F4A4", x"F44B", x"F2CE", x"F073", x"EE0C", x"EC45", x"EC55",
		x"EF01", x"F460", x"FB6C", x"02EF", x"09BB", x"0F1A", x"12BB", x"148B",
		x"151A", x"150B", x"1517", x"1549", x"1521", x"1434", x"11D2", x"0DAA",
		x"0799", x"0025", x"F858", x"F1BA", x"EDA3", x"ECC7", x"EF84", x"F4F7",
		x"FC65", x"040D", x"0AF2", x"1027", x"1352", x"14C3", x"1510", x"14B5",
		x"1415", x"133C", x"1213", x"108D", x"0E9C", x"0B83", x"06AA", x"0050",
		x"F934", x"F2C2", x"EE1C", x"EC41", x"ED2D", x"F049", x"F475", x"F86E",
		x"FB34", x"FC9C", x"FD53", x"FE62", x"00C7", x"04B0", x"09AF", x"0E76",
		x"11AC", x"1222", x"0F58", x"09F7", x"0376", x"FE0F", x"FBAB", x"FD6E",
		x"02C0", x"09A0", x"0FAA", x"12AC", x"123D", x"0FBD", x"0D29", x"0C13",
		x"0D5B", x"1008", x"126C", x"1273", x"0F09", x"081C", x"FF87", x"F712",
		x"F07F", x"EC7E", x"EB53", x"ECBD", x"F09B", x"F696", x"FDED", x"05B0",
		x"0C90", x"1196", x"13BD", x"12D0", x"0F56", x"09CF", x"037D", x"FD4F",
		x"F7D6", x"F393", x"F055", x"EE0B", x"ECC8", x"EC21", x"EBD8", x"EB7F",
		x"EB46", x"EB2E", x"EB58", x"EC06", x"ED22", x"EEC7", x"F138", x"F4B8",
		x"F963", x"FF32", x"05A9", x"0BD4", x"10B4", x"1340", x"12FC", x"0FB6",
		x"0A08", x"02D7", x"FB33", x"F468", x"EF22", x"EC3B", x"EBBA", x"EE2F",
		x"F341", x"FA5D", x"0279", x"0A6E", x"109B", x"13E7", x"13C1", x"10F1",
		x"0CF4", x"09B9", x"0863", x"0951", x"0BB9", x"0E7C", x"10E7", x"12DE",
		x"1471", x"14EB", x"137E", x"0F5C", x"089B", x"005A", x"F826", x"F144",
		x"EC79", x"E9CA", x"E927", x"EA95", x"EE1A", x"F39E", x"FAD7", x"02EC",
		x"0A9C", x"107B", x"1388", x"1357", x"1023", x"0AA7", x"0376", x"FB72",
		x"F3F1", x"EE73", x"EBC7", x"EC1A", x"EE59", x"F137", x"F3A3", x"F57D",
		x"F69D", x"F76B", x"F7B4", x"F79E", x"F715", x"F62C", x"F4DE", x"F339",
		x"F146", x"EF26", x"ED47", x"EBF3", x"EB28", x"EAFD", x"EB49", x"EBE4",
		x"ECCA", x"EDBE", x"EE88", x"EF1E", x"EF33", x"EF17", x"EEB1", x"EE1C",
		x"ED44", x"EC1F", x"EB3E", x"EB33", x"ECCB", x"F0C2", x"F73E", x"FF5E",
		x"07B4", x"0E7C", x"12CF", x"14E1", x"1559", x"1528", x"1513", x"152B",
		x"14C8", x"13CB", x"1233", x"1107", x"10F4", x"11A9", x"12C6", x"132E",
		x"11AB", x"0D45", x"0611", x"FDA7", x"F606", x"F0A3", x"ED99", x"EC3D",
		x"EBD3", x"EB9D", x"EB55", x"EAFA", x"EB1A", x"EC59", x"EF83", x"F4FA",
		x"FC7E", x"04C1", x"0C21", x"1171", x"1451", x"1540", x"154A", x"14E8",
		x"14D1", x"14D6", x"14DD", x"1452", x"130E", x"114F", x"0F3F", x"0D3B",
		x"0B41", x"0982", x"07D6", x"060B", x"03BA", x"005F", x"FBB9", x"F64E",
		x"F120", x"ED7B", x"EC2D", x"ED65", x"F134", x"F74E", x"FEE7", x"06C1",
		x"0D9A", x"1238", x"13EF", x"1274", x"0E2E", x"085F", x"0268", x"FD40",
		x"F951", x"F683", x"F48D", x"F33C", x"F220", x"F075", x"EE62", x"EC41",
		x"EB78", x"ED77", x"F295", x"F9E9", x"01FC", x"0959", x"0EE3", x"11F4",
		x"11BA", x"0DEB", x"070C", x"FECE", x"F6BF", x"F076", x"EC5C", x"EA39",
		x"E9B4", x"EAAE", x"ED33", x"F1AC", x"F85F", x"00BA", x"0933", x"0FBE",
		x"12A8", x"113B", x"0BED", x"0420", x"FB8D", x"F405", x"EE7A", x"EB5C",
		x"EA27", x"EA2B", x"EAFA", x"ECEA", x"F0CC", x"F715", x"FF2D", x"07A9",
		x"0E8B", x"1301", x"14E5", x"14F0", x"1452", x"1381", x"12E5", x"126F",
		x"124B", x"122E", x"1258", x"12F3", x"13C2", x"1498", x"14ED", x"14F0",
		x"1464", x"136C", x"121E", x"1076", x"0EA8", x"0CCB", x"0ABA", x"0866",
		x"05C6", x"0326", x"009E", x"FE76", x"FC92", x"FAED", x"F972", x"F78A",
		x"F4F2", x"F1D3", x"EE9E", x"EC6C", x"EC40", x"EEE2", x"F430", x"FB3D",
		x"02CF", x"0972", x"0DF8", x"1024", x"1031", x"0E90", x"0BFE", x"08BC",
		x"0540", x"024A", x"0112", x"0219", x"0559", x"0A05", x"0EB6", x"1205",
		x"12A4", x"0FE1", x"0A05", x"0244", x"FA23", x"F359", x"EE93", x"EC35",
		x"EC2E", x"EEA5", x"F375", x"FA56", x"027B", x"0A26", x"100D", x"12EA",
		x"12B9", x"0FF6", x"0BD4", x"0786", x"0421", x"0274", x"0273", x"0410",
		x"06D0", x"0A17", x"0D6E", x"103F", x"125B", x"13AC", x"1450", x"14AE",
		x"14D5", x"150C", x"150D", x"1493", x"12D6", x"0EE1", x"084D", x"FFD0",
		x"F71B", x"F039", x"EC31", x"EADE", x"EADF", x"EB30", x"EB64", x"EBF5",
		x"EE09", x"F275", x"F90F", x"0107", x"08BA", x"0EF0", x"12E3", x"14A7",
		x"14BD", x"13C9", x"12A1", x"11F5", x"1227", x"1326", x"1407", x"13B8",
		x"116E", x"0CD2", x"0612", x"FE3A", x"F6CD", x"F16E", x"EF7B", x"F164",
		x"F6C5", x"FE88", x"06C6", x"0DFE", x"12A5", x"147E", x"1417", x"12FF",
		x"1285", x"1302", x"141D", x"1482", x"1428", x"1371", x"1351", x"1380",
		x"135B", x"118F", x"0D50", x"06C8", x"FECB", x"F71C", x"F157", x"EE35",
		x"ED3E", x"ED9A", x"EED0", x"F0B6", x"F383", x"F6F4", x"FAB0", x"FE7B",
		x"022D", x"05A3", x"08DC", x"0B76", x"0DA0", x"0F34", x"1061", x"1100",
		x"10C2", x"0F9A", x"0D97", x"0B36", x"08A6", x"060C", x"0374", x"0162",
		x"0030", x"004C", x"01C1", x"044A", x"0771", x"0A9A", x"0D5A", x"0FA7",
		x"114A", x"1280", x"137A", x"142F", x"14C6", x"152C", x"1553", x"14EC",
		x"138A", x"1050", x"0AC7", x"034E", x"FB0B", x"F3B7", x"EE6F", x"EB95",
		x"EAEC", x"EB65", x"EC0F", x"EC34", x"EBBB", x"EB10", x"EADF", x"EB95",
		x"ECEB", x"EE8E", x"F01D", x"F1A6", x"F307", x"F486", x"F697", x"F961",
		x"FCF2", x"0142", x"0612", x"0B28", x"0FC1", x"1325", x"141C", x"1227",
		x"0D04", x"0563", x"FCF5", x"F53A", x"EFA5", x"ECE1", x"ED00", x"EFC8",
		x"F435", x"F90A", x"FD1E", x"FFD2", x"0116", x"00EE", x"FF8A", x"FCD0",
		x"F932", x"F4C5", x"F066", x"ED2E", x"EC5B", x"EEA9", x"F3D6", x"FAEE",
		x"0242", x"08BA", x"0CF9", x"0E20", x"0B8B", x"0566", x"FD56", x"F56A",
		x"EF93", x"EC8C", x"EBB2", x"EBF9", x"EC4F", x"EC86", x"ED8E", x"F0C1",
		x"F6FC", x"FF48", x"07AD", x"0D9B", x"1056", x"103C", x"0E0D", x"0A98",
		x"0693", x"02A2", x"FFAC", x"FE82", x"FFCC", x"037D", x"08C8", x"0E66",
		x"1256", x"1346", x"10E1", x"0C01", x"060C", x"002C", x"FB1C", x"F70C",
		x"F44A", x"F293", x"F1A4", x"F12F", x"F100", x"F127", x"F1C4", x"F2FD",
		x"F4B6", x"F6E7", x"F9AB", x"FCF1", x"009C", x"0433", x"0753", x"0A3F",
		x"0CC1", x"0EF3", x"10B4", x"11D7", x"1289", x"12D8", x"130E", x"1303",
		x"12C2", x"11EC", x"1049", x"0DA7", x"09D7", x"04CD", x"FEF5", x"F8B2",
		x"F2A7", x"EE11", x"EBC9", x"EC68", x"EF8B", x"F499", x"FA54", x"FFFF",
		x"0504", x"0921", x"0C4B", x"0E54", x"0F28", x"0EC9", x"0D28", x"09DC",
		x"047D", x"FDB2", x"F695", x"F0AD", x"ED21", x"EC75", x"EE2F", x"F175",
		x"F4E5", x"F7B3", x"F973", x"FA8B", x"FB8B", x"FD63", x"00E2", x"05F4",
		x"0B8D", x"1012", x"1239", x"10FF", x"0CC2", x"06E9", x"01C9", x"FF3C",
		x"004B", x"04A1", x"0A97", x"0FF3", x"12C9", x"123C", x"0E9C", x"094E",
		x"03EF", x"FF8C", x"FC6B", x"FA5B", x"F8BB", x"F6F8", x"F4D0", x"F228",
		x"EF4D", x"ECE2", x"EBCB", x"ECB6", x"EFEF", x"F582", x"FCCA", x"04C2",
		x"0C34", x"1181", x"139A", x"127D", x"0EBA", x"091C", x"0294", x"FC02",
		x"F619", x"F150", x"EDE3", x"EBC6", x"EAF4", x"EB2C", x"EBA5", x"EBDA",
		x"EB8C", x"EB63", x"EC8C", x"F008", x"F630", x"FDED", x"05CE", x"0C4F",
		x"10A7", x"12D0", x"12D6", x"10C2", x"0C71", x"05DD", x"FDE2", x"F5F1",
		x"EFCB", x"ED0F", x"EEA0", x"F446", x"FC89", x"0565", x"0CD3", x"11D6",
		x"148E", x"15CE", x"15D8", x"14B8", x"11FB", x"0D4A", x"069B", x"FE97",
		x"F698", x"F020", x"EC40", x"EAF4", x"EAFE", x"EBAB", x"ECB2", x"EE57",
		x"F0A6", x"F3C3", x"F771", x"FB58", x"FF67", x"033A", x"06AA", x"098C",
		x"0BBA", x"0CEE", x"0CE1", x"0B0D", x"0727", x"015D", x"FA6A", x"F3A0",
		x"EE9B", x"EC73", x"ED5D", x"F093", x"F4CD", x"F8F1", x"FBF0", x"FDFD",
		x"FF98", x"0125", x"02EA", x"0534", x"082D", x"0B87", x"0EE2", x"1197",
		x"135B", x"145E", x"14F8", x"1504", x"13E4", x"10E0", x"0B88", x"043B",
		x"FC1E", x"F491", x"EED6", x"EB62", x"EA0C", x"EA10", x"EA98", x"EB3C",
		x"EC0B", x"ED3C", x"EED9", x"F048", x"F0C9", x"EFE5", x"EE2A", x"EC8E",
		x"EC83", x"EF0F", x"F469", x"FC0C", x"0493", x"0C4D", x"118C", x"1351",
		x"1193", x"0CDF", x"0684", x"FFCE", x"FA28", x"F66D", x"F49E", x"F4C5",
		x"F673", x"F962", x"FD10", x"00F1", x"044B", x"0680", x"0767", x"06E5",
		x"053D", x"0295", x"FF56", x"FB96", x"F7E8", x"F4B4", x"F26B", x"F0C6",
		x"EF96", x"EEAD", x"EDA9", x"EC7A", x"EB57", x"EAA3", x"EB2C", x"ED98",
		x"F265", x"F940", x"0140", x"08FD", x"0F23", x"1329", x"1542", x"15EE",
		x"15DF", x"154F", x"144E", x"12F6", x"112A", x"0F35", x"0D86", x"0CA7",
		x"0D1D", x"0EC1", x"112B", x"1327", x"1469", x"14FD", x"155C", x"154F",
		x"1499", x"12A0", x"0ECF", x"08F5", x"0154", x"F921", x"F206", x"ED84",
		x"ECC4", x"EFCB", x"F5E5", x"FD92", x"0530", x"0BA6", x"105A", x"134B",
		x"14BF", x"151D", x"14D3", x"144A", x"134A", x"11D4", x"0FB9", x"0D24",
		x"0A0B", x"066C", x"02DA", x"FF6D", x"FC8A", x"FA05", x"F7FC", x"F66D",
		x"F5DB", x"F690", x"F85A", x"FB2F", x"FEBC", x"0273", x"05DD", x"0835",
		x"08D8", x"0729", x"02E0", x"FC59", x"F4F8", x"EF1E", x"EC8E", x"ED2D",
		x"EFD5", x"F266", x"F3B5", x"F386", x"F1C1", x"EF67", x"ECF9", x"EB55",
		x"EA63", x"EA6B", x"EB7E", x"EE4F", x"F34B", x"FA2F", x"0220", x"09E0",
		x"0FFA", x"13A5", x"1518", x"1555", x"1506", x"1491", x"13BF", x"124E",
		x"1029", x"0D7B", x"0A6F", x"073D", x"041C", x"0127", x"FE3F", x"FB80",
		x"F92D", x"F781", x"F69B", x"F680", x"F72E", x"F8C4", x"FB27", x"FDF4",
		x"0114", x"043A", x"0786", x"0A97", x"0D28", x"0F10", x"108E", x"11CC",
		x"12F0", x"13D6", x"1475", x"14DF", x"14F8", x"14BF", x"1464", x"140A",
		x"1344", x"1205", x"0FC1", x"0C26", x"06D6", x"0012", x"F887", x"F1C1",
		x"ED26", x"EB7E", x"EC93", x"EF1C", x"F1AF", x"F35E", x"F3C7", x"F307",
		x"F17D", x"EF8F", x"EDAE", x"EC4A", x"EC01", x"ED36", x"F06F", x"F5BD",
		x"FCA9", x"0432", x"0B6A", x"10C2", x"1381", x"12F8", x"0FA7", x"0A24",
		x"0359", x"FC50", x"F5B4", x"F060", x"ED4C", x"ECEE", x"EF92", x"F529",
		x"FCB1", x"04AD", x"0BA0", x"1092", x"137C", x"14D5", x"153C", x"1557",
		x"156B", x"1513", x"1438", x"1283", x"0FC6", x"0BDB", x"06C2", x"00B3",
		x"FA55", x"F46D", x"EF88", x"EC6C", x"EBE9", x"EEAB", x"F4B7", x"FD3B",
		x"065D", x"0E0D", x"12AA", x"140C", x"131E", x"1161", x"1064", x"10C7",
		x"1258", x"13AE", x"131D", x"0F97", x"0916", x"011A", x"F93E", x"F2D0",
		x"EEA6", x"EC3F", x"EB5A", x"EB0A", x"EB12", x"EAFE", x"EAE5", x"EB18",
		x"EC00", x"EE4D", x"F260", x"F864", x"0010", x"081F", x"0EAF", x"1280",
		x"1296", x"0F03", x"089A", x"00DD", x"F957", x"F359", x"EF5D", x"ECF7",
		x"EBB9", x"EB25", x"EB0E", x"EB59", x"EC1F", x"EDC9", x"F097", x"F50F",
		x"FB1A", x"0246", x"097C", x"0F5C", x"12D9", x"1398", x"1204", x"0F06",
		x"0BD3", x"0958", x"0805", x"0833", x"0980", x"0BDC", x"0EC3", x"11BC",
		x"13F5", x"144A", x"120C", x"0CEC", x"05DE", x"FDF3", x"F6B8", x"F0EF",
		x"ED36", x"EB72", x"EB46", x"EC14", x"ED9C", x"EFAD", x"F253", x"F51C",
		x"F6FB", x"F6D3", x"F47C", x"F0C9", x"ED77", x"EC5C", x"EEB5", x"F452",
		x"FBAF", x"02C5", x"0840", x"0BB9", x"0DD8", x"0F61", x"1070", x"115B",
		x"1277", x"139B", x"1457", x"13AD", x"10D4", x"0B6F", x"043C", x"FC88",
		x"F571", x"F00C", x"ECB8", x"EB1C", x"EAF8", x"EBA7", x"EC94", x"ED7F",
		x"EE72", x"EF6B", x"F082", x"F1C9", x"F345", x"F51B", x"F72D", x"F986",
		x"FC2F", x"FF79", x"036A", x"0830", x"0D01", x"1124", x"137D", x"134B",
		x"107C", x"0B1A", x"03FD", x"FC1B", x"F4C2", x"EF34", x"EC4A", x"EC0B",
		x"EE5E", x"F2ED", x"F958", x"00CE", x"0838", x"0E4B", x"1241", x"13E2",
		x"12EF", x"0F9A", x"09E3", x"02B9", x"FAE2", x"F3BF", x"EEB1", x"ECFC",
		x"EF2E", x"F471", x"FA9C", x"FF86", x"013E", x"FF3A", x"FA0F", x"F3D3",
		x"EF03", x"ED74", x"EF49", x"F2C5", x"F58D", x"F5D5", x"F380", x"F000",
		x"ED8F", x"EE42", x"F270", x"F8AD", x"FE4D", x"0111", x"FFF8", x"FBA6",
		x"F58A", x"EFEE", x"ECDB", x"EDC3", x"F2A1", x"FA27", x"02C0", x"0A80",
		x"104C", x"138A", x"13EF", x"1210", x"0E53", x"098A", x"044A", x"FF4E",
		x"FB1B", x"F7FA", x"F5E3", x"F47B", x"F34C", x"F1F9", x"F08B", x"EF14",
		x"EDC5", x"EC80", x"EB87", x"EB0B", x"EB09", x"EB57", x"EBCF", x"EC79",
		x"ED10", x"EDE5", x"EEFB", x"F0A1", x"F314", x"F697", x"FB36", x"00AF",
		x"068D", x"0C2E", x"10CE", x"137B", x"13D4", x"1102", x"0B38", x"030E",
		x"FA24", x"F273", x"EDA4", x"ECBF", x"EF23", x"F321", x"F680", x"F781",
		x"F5C9", x"F224", x"EE76", x"ECDF", x"EE9F", x"F344", x"F91E", x"FDB5",
		x"FF34", x"FD4B", x"F8D4", x"F37D", x"EF03", x"ED1F", x"EF19", x"F4EF",
		x"FD9E", x"0703", x"0EDA", x"131A", x"1372", x"10BD", x"0CB8", x"0943",
		x"07CE", x"0916", x"0C7E", x"107C", x"12DF", x"1204", x"0DEC", x"07F9",
		x"01FC", x"FDB0", x"FBE9", x"FCB9", x"FFA5", x"03DA", x"0856", x"0C6D",
		x"0F88", x"1181", x"12D0", x"13AC", x"1465", x"14E3", x"1528", x"1502",
		x"144C", x"126F", x"0EBF", x"0943", x"0262", x"FB04", x"F43C", x"EF25",
		x"EC48", x"EBD2", x"ED0F", x"EF5B", x"F202", x"F434", x"F5E3", x"F73C",
		x"F8A7", x"FA7C", x"FD05", x"000D", x"03BD", x"07E8", x"0BE6", x"0F23",
		x"111D", x"11AB", x"1028", x"0C2B", x"057B", x"FD25", x"F504", x"EF3D",
		x"EC7A", x"EBCF", x"EBD9", x"EBC6", x"EBEC", x"ED11", x"F07E", x"F677",
		x"FE76", x"0677", x"0C66", x"0F06", x"0DD8", x"09BD", x"036C", x"FBEF",
		x"F49F", x"EF14", x"ECEF", x"EECC", x"F48A", x"FCCD", x"0578", x"0CBF",
		x"1193", x"13F1", x"1472", x"13EB", x"1314", x"12C8", x"1330", x"141B",
		x"14D3", x"14E4", x"1465", x"13D2", x"1379", x"1375", x"13E3", x"1471",
		x"14CE", x"149D", x"13FE", x"1344", x"12C6", x"12A6", x"12EA", x"1370",
		x"140D", x"14B2", x"14E7", x"145B", x"12A2", x"0F36", x"09F8", x"032C",
		x"FBBB", x"F4CF", x"EF81", x"EC8C", x"EBF2", x"ED52", x"EFD6", x"F312",
		x"F66F", x"F95A", x"FBED", x"FD92", x"FE40", x"FDF6", x"FCB9", x"FAD0",
		x"F88E", x"F623", x"F3CA", x"F19E", x"EFC2", x"EE76", x"EDEE", x"EE0E",
		x"EE8A", x"EF68", x"F0CE", x"F353", x"F6F4", x"FC16", x"021B", x"08A5",
		x"0E7C", x"125A", x"12FA", x"1046", x"0BA2", x"071D", x"04A0", x"0550",
		x"08D7", x"0DAA", x"11B8", x"12ED", x"10C9", x"0BA6", x"04FC", x"FE1F",
		x"F82C", x"F422", x"F1BC", x"F077", x"EFCE", x"EF56", x"EF11", x"EF10",
		x"EF60", x"EFC6", x"F074", x"F1AB", x"F3CC", x"F6EF", x"FB51", x"00EF",
		x"071C", x"0D0D", x"1171", x"131A", x"11C0", x"0DBC", x"0894", x"03ED",
		x"0132", x"00E4", x"02BB", x"0609", x"09E5", x"0D93", x"1009", x"10FC",
		x"0FF1", x"0C3F", x"05F1", x"FDFC", x"F616", x"F00F", x"ECCC", x"EBE7",
		x"EC4F", x"ECF7", x"ECFC", x"EC5A", x"EBAD", x"EB74", x"EBBE", x"EBEF",
		x"EBA7", x"EB27", x"EB72", x"ED9B", x"F23E", x"F912", x"00FC", x"087F",
		x"0E21", x"1178", x"12D1", x"12A3", x"117D", x"0F6A", x"0C9C", x"091B",
		x"0557", x"01BD", x"FE5C", x"FB80", x"F90D", x"F719", x"F55A", x"F3C4",
		x"F1FA", x"F019", x"EE4F", x"ECC9", x"EBB4", x"EAF6", x"EA8A", x"EA7A",
		x"EB07", x"EBFE", x"ED27", x"EE58", x"EFE8", x"F1B8", x"F3D9", x"F612",
		x"F87A", x"FB19", x"FDAD", x"0009", x"01D9", x"0343", x"048D", x"0636",
		x"08A7", x"0BD6", x"0F69", x"1244", x"1365", x"11CE", x"0D46", x"0668",
		x"FEC8", x"F80B", x"F3AA", x"F22C", x"F3B9", x"F7E3", x"FE25", x"0573",
		x"0C61", x"113F", x"12A1", x"102F", x"0AA5", x"0386", x"FC31", x"F58A",
		x"F04D", x"ED16", x"EC43", x"EE45", x"F2BD", x"F907", x"0030", x"075F",
		x"0DA2", x"122B", x"1427", x"1329", x"0F1D", x"087C", x"0015", x"F7A7",
		x"F0D9", x"ECAF", x"EB57", x"EBDF", x"ECF9", x"EDAF", x"ED83", x"ECCE",
		x"EBE6", x"EB5C", x"EB45", x"EB57", x"EB3D", x"EAF9", x"EB2D", x"ECB6",
		x"F09E", x"F6F3", x"FF3E", x"07E3", x"0F16", x"1350", x"142A", x"11F1",
		x"0D62", x"0734", x"0015", x"F8D5", x"F28A", x"EE27", x"EC5C", x"EDA1",
		x"F1D3", x"F83D", x"FFAC", x"06D0", x"0CD5", x"10F0", x"1396", x"149B",
		x"149D", x"13E1", x"12D9", x"1202", x"1196", x"117E", x"11A9", x"11E0",
		x"1215", x"1274", x"131E", x"1404", x"14BA", x"14CC", x"135B", x"0F93",
		x"0930", x"00E4", x"F856", x"F189", x"ED43", x"EB3F", x"EA7D", x"EA55",
		x"EABF", x"EC6D", x"F027", x"F683", x"FED1", x"0782", x"0E88", x"1265",
		x"1249", x"0E94", x"082D", x"0099", x"F913", x"F2E5", x"EEBA", x"EC8B",
		x"EBFD", x"EC91", x"EDE6", x"F021", x"F336", x"F689", x"F8CE", x"F917",
		x"F6FC", x"F330", x"EF42", x"ED26", x"EE56", x"F30D", x"F98C", x"FFB2",
		x"03CA", x"04D4", x"0345", x"FFE3", x"FBBC", x"F7C2", x"F499", x"F2F2",
		x"F355", x"F638", x"FB65", x"0238", x"097D", x"0F85", x"1311", x"13AB",
		x"1176", x"0D60", x"08AF", x"0461", x"010E", x"FEB1", x"FD13", x"FC0A",
		x"FBB5", x"FBDC", x"FC9A", x"FDFC", x"FFF9", x"0247", x"04E8", x"07DB",
		x"0AC7", x"0D7A", x"0FBC", x"117D", x"12E7", x"13EE", x"14A4", x"1520",
		x"153A", x"1502", x"1490", x"13FD", x"133D", x"1242", x"10F0", x"0F1E",
		x"0C73", x"08BB", x"03FD", x"FE3A", x"F7E7", x"F20A", x"EDC2", x"EC23",
		x"ED5A", x"F0CF", x"F5E0", x"FB90", x"0153", x"063C", x"09E6", x"0C13",
		x"0CF2", x"0CB4", x"0B54", x"0891", x"0445", x"FE8B", x"F82D", x"F22C",
		x"EDD7", x"EC6C", x"EEA4", x"F421", x"FB7F", x"0328", x"0A0E", x"0F8E",
		x"132F", x"1462", x"12B9", x"0E19", x"06D9", x"FE0A", x"F566", x"EEC3",
		x"EB7A", x"EB59", x"ECF1", x"EE6D", x"EEB2", x"EDB3", x"EC77", x"ECB0",
		x"F003", x"F675", x"FEC3", x"06B2", x"0CCC", x"108F", x"12A8", x"1370",
		x"13AF", x"13D9", x"143B", x"14BE", x"1481", x"124F", x"0D2D", x"05A6",
		x"FD0B", x"F545", x"EF95", x"EC15", x"EA60", x"EA1E", x"EB90", x"EF08",
		x"F4CD", x"FC5B", x"04B0", x"0C56", x"11C0", x"143C", x"1499", x"13E6",
		x"135C", x"131C", x"12D0", x"11EB", x"0FE9", x"0C36", x"0654", x"FED3",
		x"F6E9", x"F07F", x"ED15", x"ECD5", x"EE50", x"EFA1", x"EF91", x"EE12",
		x"EC59", x"EC12", x"EECA", x"F45A", x"FBD9", x"03C7", x"0AA7", x"0FCC",
		x"12F3", x"14A9", x"152F", x"1549", x"1560", x"157B", x"154D", x"13BC",
		x"1002", x"09B3", x"01E6", x"F9DD", x"F2EA", x"EE01", x"EB5A", x"EAEF",
		x"ECAF", x"F0A1", x"F6AC", x"FE80", x"06BD", x"0DF9", x"12DE", x"14BF",
		x"13D9", x"1171", x"0E97", x"0C03", x"0A26", x"0942", x"09BC", x"0BC2",
		x"0EBE", x"11B9", x"1335", x"122D", x"0E26", x"07F0", x"0121", x"FB68",
		x"F7CD", x"F682", x"F739", x"F930", x"FC34", x"FFD9", x"03EB", x"080E",
		x"0BE2", x"0F28", x"118E", x"1351", x"147A", x"1505", x"1536", x"1548",
		x"1509", x"13DB", x"10C7", x"0B6C", x"041A", x"FC15", x"F4AA", x"EF1B",
		x"EBC4", x"EA66", x"EA1D", x"EA6B", x"EAF3", x"EC38", x"EE35", x"F0E7",
		x"F3E7", x"F6E3", x"F974", x"FB5C", x"FCA3", x"FD96", x"FEEC", x"017F",
		x"0572", x"0A45", x"0EE8", x"1247", x"135D", x"113A", x"0C28", x"052C",
		x"FE61", x"F97B", x"F6ED", x"F6B9", x"F84B", x"FB36", x"FEC6", x"026A",
		x"05BD", x"0844", x"09CB", x"0A55", x"09B5", x"0841", x"064B", x"03B4",
		x"0036", x"FBA8", x"F662", x"F141", x"ED91", x"ECB2", x"EF3A", x"F4C6",
		x"FBCE", x"021A", x"05B9", x"058B", x"01C0", x"FB76", x"F4B2", x"EF79",
		x"ED18", x"EDEF", x"F0B1", x"F3E0", x"F5E7", x"F626", x"F4EC", x"F289",
		x"EFD7", x"ED6A", x"EBB4", x"EAE4", x"EAE8", x"EBC3", x"ED21", x"EEEB",
		x"F0DB", x"F274", x"F328", x"F27C", x"F085", x"EE20", x"EC86", x"ED2F",
		x"F0DC", x"F71D", x"FEB8", x"05A8", x"0A23", x"0BB9", x"0AB7", x"0816",
		x"042D", x"FF94", x"FB43", x"F84B", x"F731", x"F818", x"FAC2", x"FE63",
		x"02BD", x"06A6", x"09BF", x"0B3C", x"0AC6", x"07DE", x"026F", x"FB3F",
		x"F40D", x"EECF", x"EC6C", x"ECEB", x"EF15", x"F160", x"F29C", x"F257",
		x"F0CA", x"EEC4", x"ECE7", x"EB98", x"EABF", x"EA68", x"EA61", x"EAA6",
		x"EB1C", x"EBCE", x"ECBD", x"EE29", x"EFE3", x"F1EF", x"F476", x"F778",
		x"FACB", x"FE25", x"0144", x"03DD", x"05DC", x"06F6", x"06EC", x"05DB",
		x"03AC", x"00F2", x"FDB5", x"FA55", x"F75F", x"F553", x"F47F", x"F4B8",
		x"F5BB", x"F743", x"F965", x"FC06", x"FF0B", x"025D", x"05FE", x"0993",
		x"0CE3", x"0FB2", x"11D5", x"1360", x"144A", x"14BC", x"14E3", x"1415",
		x"11CC", x"0D4E", x"06D7", x"FF13", x"F780", x"F13F", x"ECFA", x"EB34",
		x"EB8B", x"ED52", x"EF98", x"F18C", x"F319", x"F45D", x"F5D3", x"F791",
		x"F995", x"FB7A", x"FD4C", x"FEF1", x"00F9", x"0388", x"06DF", x"0AEA",
		x"0F0E", x"1248", x"13E2", x"1344", x"0FFF", x"0A79", x"0358", x"FBE8",
		x"F561", x"F08E", x"ED57", x"EB95", x"EADC", x"EAD9", x"EAFB", x"EAEA",
		x"EAE3", x"EB1C", x"EC56", x"EF11", x"F39C", x"F9F6", x"01A4", x"0977",
		x"0FD9", x"12F5", x"11E5", x"0C9E", x"04C2", x"FC5B", x"F52A", x"EFED",
		x"ECBF", x"EBBA", x"ED48", x"F19B", x"F847", x"0043", x"07FD", x"0E74",
		x"12D2", x"1555", x"15EB", x"14F0", x"1230", x"0D4B", x"0623", x"FD60",
		x"F4D9", x"EE68", x"EB06", x"EA47", x"EABF", x"EB50", x"EB70", x"EB97",
		x"EC47", x"EE17", x"F173", x"F6DD", x"FE15", x"060F", x"0D24", x"11CF",
		x"1396", x"1321", x"11B6", x"1030", x"0F92", x"1005", x"113E", x"12C7",
		x"1433", x"14EC", x"14DB", x"142F", x"1317", x"120F", x"113A", x"1092",
		x"0F82", x"0DAF", x"0A87", x"05B4", x"FF3D", x"F7F6", x"F170", x"ED57",
		x"ECAC", x"EF01", x"F287", x"F524", x"F56A", x"F346", x"EFC7", x"ED0A",
		x"ECF5", x"F02C", x"F670", x"FDE8", x"04E1", x"0A17", x"0D48", x"0EC1",
		x"0F32", x"0F99", x"1074", x"1208", x"1379", x"13A8", x"116A", x"0C1E",
		x"0487", x"FC2A", x"F4BE", x"EF6E", x"ECD9", x"ED32", x"F069", x"F60F",
		x"FD6D", x"0557", x"0C94", x"11EE", x"14B6", x"154F", x"14E0", x"149C",
		x"147A", x"13E3", x"128A", x"10E7", x"102A", x"10D0", x"1233", x"12D5",
		x"1151", x"0D03", x"0688", x"FEF2", x"F81C", x"F3C8", x"F319", x"F64B",
		x"FC7A", x"0441", x"0BAF", x"1104", x"1388", x"1309", x"1031", x"0C27",
		x"07D5", x"0420", x"014D", x"FF1B", x"FDC4", x"FD12", x"FD1C", x"FE3F",
		x"0078", x"0378", x"0699", x"098B", x"0BDF", x"0DA5", x"0EC6", x"0F30",
		x"0E9C", x"0D51", x"0B77", x"093A", x"0685", x"0358", x"FF9D", x"FBA6",
		x"F7A0", x"F3FE", x"F103", x"EEAF", x"ED0F", x"EBF8", x"EBA3", x"EC87",
		x"EF64", x"F478", x"FBAE", x"03A8", x"0B0C", x"109A", x"13ED", x"1521",
		x"14F7", x"148F", x"1492", x"1501", x"1523", x"14AE", x"13B0", x"1290",
		x"11AE", x"112A", x"1145", x"1210", x"132F", x"1460", x"1503", x"14B3",
		x"12DB", x"0F2A", x"09CF", x"034C", x"FC4B", x"F57D", x"EFE3", x"EC7D",
		x"EB9B", x"ECD9", x"EF6F", x"F28F", x"F5B3", x"F82B", x"F9E4", x"FAE1",
		x"FB69", x"FB5E", x"FA87", x"F8F7", x"F6ED", x"F4EC", x"F307", x"F121",
		x"EF39", x"ED67", x"EC06", x"EB6B", x"EBA4", x"ECAC", x"EE0E", x"EF73",
		x"EFCE", x"EEE6", x"ED5B", x"ECB2", x"EE2B", x"F24C", x"F8C5", x"006C",
		x"078A", x"0C7C", x"0E47", x"0C84", x"07E2", x"0156", x"F9E9", x"F316",
		x"EE48", x"EC95", x"EE23", x"F1E0", x"F655", x"FA79", x"FDF3", x"0081",
		x"01DD", x"01AA", x"FFE3", x"FC85", x"F7F1", x"F2E5", x"EEA4", x"ECAA",
		x"EDD0", x"F198", x"F739", x"FD55", x"0312", x"0805", x"0BC0", x"0E83",
		x"1031", x"1129", x"114E", x"10CD", x"0F8D", x"0D6A", x"0AA5", x"075B",
		x"03F5", x"012B", x"FFBD", x"005C", x"0341", x"0806", x"0D64", x"11CB",
		x"138E", x"11D7", x"0DA9", x"0885", x"03EB", x"0120", x"0075", x"01B5",
		x"0459", x"07E4", x"0BE6", x"0F97", x"12A0", x"1440", x"13A5", x"10A1",
		x"0B43", x"0461", x"FD11", x"F620", x"F090", x"ECBA", x"EAE7", x"EAB4",
		x"EB73", x"EC52", x"ECE6", x"ED37", x"ED1F", x"ECCF", x"EC34", x"EB8A",
		x"EB36", x"EB01", x"EB06", x"EB58", x"EBC9", x"EC6D", x"ECCC", x"ECC4",
		x"EC3B", x"EB8E", x"EB32", x"EB5D", x"EC5E", x"EE92", x"F1F5", x"F6C8",
		x"FCBA", x"0366", x"0A29", x"0FDA", x"132B", x"1362", x"1052", x"0A8F",
		x"0326", x"FB43", x"F419", x"EEBA", x"EB9C", x"EAF8", x"EC53", x"EEEF",
		x"F22E", x"F597", x"F897", x"FB1E", x"FCBE", x"FDA6", x"FDC4", x"FD5D",
		x"FC8F", x"FB77", x"FA50", x"F8BB", x"F698", x"F3CD", x"F04E", x"ED4A",
		x"EC1A", x"EE0E", x"F344", x"FABC", x"02DE", x"09E6", x"0ED6", x"10CD",
		x"0F2F", x"0A0A", x"0256", x"F9CE", x"F270", x"ED7F", x"EB19", x"EA54",
		x"EA74", x"EB19", x"ECE8", x"F0A9", x"F714", x"FF89", x"0829", x"0EF9",
		x"1287", x"1343", x"11DE", x"0F04", x"0B2F", x"06F4", x"036F", x"01B1",
		x"0277", x"05E1", x"0B16", x"102D", x"12F3", x"1243", x"0E51", x"08E0",
		x"03F2", x"00E1", x"0040", x"01B1", x"0483", x"07D5", x"0B37", x"0E1E",
		x"1024", x"113E", x"113F", x"106D", x"0EA8", x"0C55", x"0970", x"0629",
		x"02A0", x"FEEB", x"FB60", x"F819", x"F53C", x"F2B6", x"F0AB", x"EF00",
		x"EDEB", x"ED66", x"ED63", x"EDB9", x"EEBB", x"F06F", x"F2D2", x"F5A7",
		x"F8AE", x"FBCE", x"FEFA", x"01E1", x"0488", x"06BB", x"08BF", x"0A74",
		x"0C2B", x"0E12", x"102F", x"1241", x"13D1", x"14A9", x"14C8", x"147D",
		x"1438", x"1432", x"1493", x"14B8", x"1404", x"11C9", x"0D68", x"06E1",
		x"FEEC", x"F70A", x"F0AD", x"EC9E", x"EACB", x"EA8E", x"EAD6", x"EB58",
		x"EBEE", x"EC92", x"ED66", x"EF50", x"F2C6", x"F847", x"FF47", x"06DC",
		x"0D82", x"1218", x"139D", x"1187", x"0C77", x"0592", x"FE17", x"F6F6",
		x"F141", x"ED76", x"EC1A", x"ECE5", x"EF67", x"F2F1", x"F6FA", x"FB08",
		x"FE58", x"00AE", x"01D1", x"0183", x"FFBE", x"FC6D", x"F7F1", x"F2F8",
		x"EEC7", x"ECA5", x"ED90", x"F1DA", x"F8F8", x"015C", x"0941", x"0F48",
		x"1315", x"1484", x"13D6", x"1098", x"0ACA", x"0300", x"FAA0", x"F349",
		x"EE83", x"ED4A", x"EF40", x"F2F0", x"F64A", x"F76F", x"F5CF", x"F23A",
		x"EE8A", x"EC8A", x"EDAF", x"F1C7", x"F786", x"FD69", x"01E8", x"0490",
		x"0546", x"0419", x"0153", x"FD40", x"F885", x"F399", x"EF85", x"ED00",
		x"ED2D", x"F060", x"F633", x"FD64", x"0464", x"098E", x"0BF3", x"0B24",
		x"0764", x"0156", x"FA45", x"F39D", x"EED3", x"ECEE", x"EE13", x"F180",
		x"F5B2", x"F93E", x"FB71", x"FCA6", x"FD93", x"FEF5", x"00DF", x"03C0",
		x"0740", x"0B05", x"0E86", x"1144", x"131B", x"1405", x"1406", x"1317",
		x"10CF", x"0CBD", x"06B0", x"FF3D", x"F7AC", x"F13B", x"ED1F", x"EB80",
		x"EC4F", x"EED1", x"F262", x"F61B", x"F944", x"FB40", x"FBB6", x"FA6D",
		x"F78F", x"F384", x"EF7B", x"ED4D", x"EE36", x"F27B", x"F88A", x"FE4B",
		x"0156", x"0077", x"FC08", x"F5A3", x"F017", x"ED88", x"EE81", x"F1DB",
		x"F5D1", x"F893", x"F916", x"F781", x"F467", x"F103", x"EE19", x"EC52",
		x"EB92", x"EC53", x"EEE6", x"F39A", x"FA51", x"0228", x"09EA", x"1025",
		x"13C7", x"14AC", x"13AF", x"11B3", x"0FCD", x"0E24", x"0CDB", x"0BAD",
		x"0A10", x"07CF", x"0511", x"020C", x"FEC9", x"FB6C", x"F832", x"F58F",
		x"F3C3", x"F2CF", x"F2DF", x"F3E3", x"F5AC", x"F80C", x"FACF", x"FDBE",
		x"00A5", x"02FA", x"0475", x"04FF", x"04AB", x"035F", x"013F", x"FE3A",
		x"FAA6", x"F6C1", x"F2F5", x"EF7C", x"ECE0", x"EC01", x"ED0F", x"F0A4",
		x"F678", x"FE1C", x"065A", x"0D9A", x"1253", x"138B", x"1123", x"0C0E",
		x"05A0", x"FF24", x"F996", x"F5A3", x"F394", x"F34B", x"F493", x"F6E3",
		x"FA38", x"FE1A", x"021F", x"05DA", x"0906", x"0B73", x"0D1E", x"0E32",
		x"0F06", x"1019", x"11A5", x"1366", x"145B", x"12E5", x"0E47", x"06F0",
		x"FE70", x"F6C2", x"F0C8", x"ED01", x"EB7D", x"EC83", x"F026", x"F635",
		x"FE01", x"0661", x"0DAB", x"12C3", x"1549", x"15D1", x"1587", x"14F5",
		x"140B", x"123F", x"0FFA", x"0E37", x"0DC0", x"0F0F", x"1130", x"12A8",
		x"11DB", x"0E26", x"07BD", x"0018", x"F990", x"F651", x"F77A", x"FC8E",
		x"03D2", x"0B2E", x"1084", x"131E", x"12CD", x"10CA", x"0E8D", x"0D7F",
		x"0E11", x"0FDB", x"1219", x"13DF", x"150C", x"1584", x"1599", x"156A",
		x"1515", x"1483", x"136E", x"11C9", x"0FDF", x"0E1A", x"0D11", x"0D26",
		x"0E36", x"0FBB", x"1137", x"128B", x"13A3", x"146F", x"14D2", x"14AD",
		x"13E2", x"129F", x"10ED", x"0F19", x"0D1E", x"0B6F", x"0A65", x"0A65",
		x"0B4B", x"0CDF", x"0EFB", x"114A", x"1352", x"14BB", x"1550", x"1560",
		x"150B", x"148E", x"13A5", x"125D", x"10AA", x"0EC6", x"0CEE", x"0B80",
		x"0AA3", x"0A8E", x"0B52", x"0CEF", x"0F07", x"1124", x"1303", x"141F",
		x"13FB", x"1235", x"0E5A", x"08A0", x"0188", x"F9F5", x"F32D", x"EE48",
		x"EBB5", x"EB30", x"EC0E", x"ED73", x"EEF9", x"F044", x"F188", x"F2A3",
		x"F3E6", x"F571", x"F776", x"F9F6", x"FCE3", x"FFF3", x"0328", x"0613",
		x"0896", x"0AA1", x"0C6E", x"0DEA", x"0F0A", x"0FF7", x"10F7", x"1266",
		x"13FF", x"1489", x"12D8", x"0E18", x"06E7", x"FE97", x"F6EB", x"F13D",
		x"ED8F", x"EBC8", x"EB7A", x"EC83", x"EF1C", x"F3A5", x"FA7A", x"02B8",
		x"0ACC", x"1091", x"125C", x"0FB8", x"098F", x"0189", x"F987", x"F30D",
		x"EEBA", x"EC71", x"EBBD", x"EC2E", x"EDD4", x"F12C", x"F6C2", x"FE77",
		x"0720", x"0E9A", x"12DF", x"12C9", x"0E76", x"0744", x"FF16", x"F760",
		x"F155", x"ED7E", x"EBB3", x"EB05", x"EAFA", x"EB4E", x"EC1B", x"EDA9",
		x"EFC7", x"F1ED", x"F309", x"F2B7", x"F103", x"EEAE", x"ED24", x"EDE6",
		x"F195", x"F82C", x"003B", x"07CC", x"0D2F", x"104C", x"11D1", x"1293",
		x"1348", x"141B", x"14D1", x"150D", x"1448", x"11CC", x"0D3F", x"06B8",
		x"FF1D", x"F799", x"F13E", x"ED2A", x"EB56", x"EB8A", x"ED0B", x"EF07",
		x"F0CA", x"F25A", x"F39F", x"F4AF", x"F55E", x"F564", x"F4C1", x"F37A",
		x"F1F0", x"F03F", x"EE82", x"ECEA", x"EBAA", x"EB85", x"ECC3", x"EFDE",
		x"F507", x"FBD3", x"039F", x"0B0A", x"10CD", x"13CB", x"13C1", x"10D2",
		x"0BA1", x"050D", x"FDD5", x"F6C0", x"F0F4", x"ED39", x"EC44", x"EE68",
		x"F35C", x"FA48", x"01AF", x"08AF", x"0E39", x"1225", x"145A", x"14EC",
		x"1413", x"1225", x"0FA8", x"0D55", x"0C25", x"0C7C", x"0E62", x"10C0",
		x"1258", x"11D8", x"0E71", x"0870", x"0117", x"FA6A", x"F65F", x"F65D",
		x"FA98", x"01BC", x"0983", x"0F84", x"12B4", x"133B", x"1273", x"11A0",
		x"11C2", x"12AD", x"1388", x"1269", x"0E1C", x"06CD", x"FDB4", x"F50D",
		x"EF07", x"EC96", x"EDCF", x"F209", x"F808", x"FE7A", x"046C", x"08F2",
		x"0BEB", x"0D36", x"0CE2", x"0B30", x"084B", x"0499", x"0074", x"FC6E",
		x"F882", x"F51E", x"F256", x"F019", x"EE7D", x"ED5C", x"EC9A", x"EC2B",
		x"EC02", x"EBF5", x"EBE6", x"EC28", x"ECA5", x"EDD4", x"EFF2", x"F379",
		x"F866", x"FE75", x"0548", x"0BC0", x"10B5", x"1378", x"139E", x"1159",
		x"0D41", x"07E0", x"01EA", x"FC34", x"F781", x"F41A", x"F1C6", x"F0CD",
		x"F140", x"F375", x"F7DD", x"FE2D", x"056E", x"0C23", x"111F", x"13A1",
		x"13F1", x"12B0", x"10C6", x"0F2D", x"0E90", x"0F36", x"10C8", x"12C1",
		x"1455", x"14A6", x"12AB", x"0E17", x"06FD", x"FE9C", x"F6C1", x"F0C8",
		x"ED19", x"EB3A", x"EA88", x"EAAA", x"EBD6", x"EED0", x"F426", x"FBA0",
		x"0446", x"0C3C", x"11E5", x"14D4", x"1566", x"14DA", x"13FB", x"1351",
		x"12B4", x"11F7", x"10FC", x"0F82", x"0DDE", x"0C05", x"0A2C", x"0847",
		x"0638", x"0385", x"FFC1", x"FAEA", x"F57D", x"F09D", x"ED3F", x"EC65",
		x"EE37", x"F288", x"F890", x"FF09", x"0541", x"0A49", x"0E10", x"10B6",
		x"127D", x"1395", x"141C", x"13C7", x"1235", x"0E64", x"0813", x"0013",
		x"F81C", x"F1AB", x"ED68", x"EB16", x"EA48", x"EAAA", x"ECA3", x"F093",
		x"F6C5", x"FEE5", x"076D", x"0EB8", x"131B", x"1359", x"0F81", x"08A2",
		x"004B", x"F823", x"F17D", x"ECFF", x"EAAB", x"EA0C", x"EABF", x"EC69",
		x"EFC6", x"F55C", x"FD41", x"05E9", x"0D82", x"12AA", x"153B", x"15E7",
		x"15A5", x"14FD", x"1456", x"13BF", x"131F", x"1209", x"1049", x"0DE7",
		x"0B27", x"084B", x"056E", x"02BC", x"00A0", x"FF46", x"FF00", x"FFB5",
		x"0133", x"035D", x"05D9", x"08C4", x"0BBC", x"0E88", x"10C5", x"1235",
		x"133A", x"13EF", x"14A9", x"1506", x"152C", x"14C2", x"1377", x"1065",
		x"0AD0", x"02F2", x"FA50", x"F2DE", x"EDCD", x"EB30", x"EA4F", x"EA2B",
		x"EACD", x"EC9F", x"F000", x"F588", x"FCFE", x"0536", x"0C64", x"1159",
		x"13B3", x"1429", x"138E", x"122E", x"0FDC", x"0C7D", x"07F6", x"028A",
		x"FCB2", x"F6DB", x"F1B9", x"EE05", x"EC52", x"ED32", x"F0E3", x"F71F",
		x"FF28", x"07A2", x"0ED3", x"1331", x"13FC", x"1192", x"0D31", x"0892",
		x"04FB", x"035C", x"03D2", x"05F7", x"0901", x"0C42", x"0F48", x"118A",
		x"12A7", x"127F", x"115C", x"0F2F", x"0C42", x"0906", x"05F9", x"03BC",
		x"0323", x"045C", x"078B", x"0BFA", x"1032", x"12E5", x"12CF", x"0F96",
		x"0964", x"0170", x"F91F", x"F213", x"EDD7", x"ECA0", x"EEA9", x"F2E4",
		x"F7FA", x"FC25", x"FE8A", x"FEDA", x"FD40", x"FA7A", x"F72C", x"F40F",
		x"F183", x"EF9B", x"EE67", x"EE60", x"EFA1", x"F229", x"F56E", x"F8DD",
		x"FBF3", x"FE37", x"FF2C", x"FE7E", x"FC25", x"F8A6", x"F4D8", x"F195",
		x"EF4B", x"EE1D", x"EE40", x"F049", x"F4E1", x"FBA7", x"03BA", x"0B4F",
		x"10EA", x"13E2", x"1484", x"13D7", x"131A", x"1321", x"13B5", x"1433",
		x"1433", x"13CC", x"132F", x"12BE", x"12D5", x"134E", x"142F", x"14D4",
		x"1522", x"14BE", x"13FD", x"1356", x"1300", x"1347", x"13F5", x"1490",
		x"14ED", x"14D0", x"1456", x"1346", x"1185", x"0F1D", x"0C66", x"09A9",
		x"070E", x"04B8", x"02C6", x"0175", x"00E3", x"0128", x"0236", x"03DA",
		x"05CF", x"083C", x"0AFB", x"0DBB", x"102D", x"1242", x"13E2", x"1509",
		x"158E", x"1561", x"14F6", x"1472", x"142D", x"141F", x"1427", x"1437",
		x"1469", x"14AE", x"1505", x"14D2", x"1397", x"10DD", x"0C52", x"060F",
		x"FEA6", x"F73F", x"F107", x"ED43", x"EC11", x"ED19", x"EF72", x"F21B",
		x"F497", x"F6A7", x"F878", x"FA36", x"FC9A", x"FFD7", x"0426", x"0959",
		x"0E73", x"1243", x"1359", x"113A", x"0C38", x"05CB", x"FFAA", x"FAD6",
		x"F78D", x"F592", x"F45A", x"F387", x"F270", x"F079", x"EE17", x"EC6B",
		x"ED10", x"F0C5", x"F726", x"FEEB", x"0668", x"0C81", x"1078", x"11DF",
		x"1097", x"0CCF", x"06DC", x"FF5D", x"F77B", x"F0F3", x"ED68", x"EDB7",
		x"F16A", x"F76B", x"FE6F", x"05C8", x"0C80", x"11A8", x"145F", x"144D",
		x"119F", x"0C90", x"05EF", x"FE7B", x"F752", x"F14C", x"ED54", x"EC06",
		x"EDB2", x"F212", x"F89B", x"0033", x"0790", x"0DD4", x"1250", x"148C",
		x"1497", x"12D8", x"0FCA", x"0C41", x"08F7", x"0661", x"04E8", x"04A0",
		x"05BD", x"0837", x"0BF3", x"0FE0", x"12D4", x"133D", x"1060", x"0AB5",
		x"0355", x"FB4F", x"F414", x"EECC", x"EC25", x"EC80", x"EF82", x"F484",
		x"FAFF", x"0234", x"0917", x"0EBD", x"1256", x"13AF", x"1293", x"0F1F",
		x"0920", x"013A", x"F8F4", x"F1E7", x"EDA3", x"ECAD", x"EEDF", x"F33E",
		x"F881", x"FD7E", x"0138", x"03BD", x"04CC", x"0470", x"02B6", x"FF8A",
		x"FB2D", x"F601", x"F0EB", x"ED65", x"EC6E", x"EEA6", x"F398", x"FA23",
		x"00FC", x"06CD", x"0A75", x"0B5A", x"0943", x"047C", x"FDFB", x"F6FC",
		x"F111", x"EDF0", x"EEA3", x"F308", x"FA27", x"023F", x"09ED", x"0FCD",
		x"138C", x"14C8", x"13E9", x"1125", x"0CEF", x"0820", x"0357", x"FF47",
		x"FC31", x"FA66", x"FA63", x"FC24", x"FFCB", x"04F8", x"0AC1", x"101F",
		x"1378", x"1422", x"11DE", x"0D36", x"073D", x"0100", x"FB49", x"F6C1",
		x"F3D8", x"F24D", x"F1E6", x"F265", x"F427", x"F754", x"FC24", x"0221",
		x"08B4", x"0EAD", x"12BF", x"138E", x"10A5", x"0A5A", x"01E1", x"F936",
		x"F219", x"ED8F", x"EBE2", x"EC63", x"EE1B", x"EFDE", x"F129", x"F169",
		x"F0AB", x"EF22", x"ED40", x"EBB1", x"EB0D", x"EBFE", x"EEDB", x"F3BC",
		x"FA58", x"01D5", x"0921", x"0F24", x"1316", x"14BF", x"147A", x"135D",
		x"1208", x"10F3", x"0FD0", x"0E8B", x"0C96", x"098A", x"050B", x"FF07",
		x"F83A", x"F1F0", x"EDDE", x"ED0E", x"EF3B", x"F2C7", x"F5B7", x"F6CB",
		x"F60C", x"F3D1", x"F10F", x"EE96", x"ECD1", x"EBD9", x"EBBE", x"EC81",
		x"EEAF", x"F2E2", x"F936", x"0107", x"0929", x"0FB6", x"1344", x"1332",
		x"0FE9", x"0A64", x"03B7", x"FC92", x"F5F9", x"F086", x"ECF8", x"EC19",
		x"EE3F", x"F35C", x"FA84", x"028A", x"09EB", x"0F8E", x"12F5", x"144D",
		x"1449", x"136F", x"1236", x"10A9", x"0EE1", x"0D14", x"0B45", x"0998",
		x"07EB", x"0657", x"04D1", x"034B", x"01AB", x"FF96", x"FC9B", x"F883",
		x"F3D9", x"EFAC", x"ED70", x"EDD7", x"F138", x"F706", x"FDD8", x"03C9",
		x"0770", x"07F5", x"0569", x"008A", x"FA1F", x"F394", x"EE93", x"ECF9",
		x"EF96", x"F5FB", x"FED0", x"080C", x"0F51", x"1345", x"13EB", x"1282",
		x"10E8", x"1063", x"1151", x"12DB", x"139A", x"11AA", x"0C7B", x"04CA",
		x"FCF9", x"F7D5", x"F6FE", x"FAC4", x"01A2", x"095B", x"0F73", x"125D",
		x"121F", x"0FD3", x"0D7B", x"0C88", x"0D6F", x"0FB2", x"1227", x"13E7",
		x"14B0", x"14F6", x"14CF", x"1407", x"11B1", x"0D01", x"063E", x"FE48",
		x"F68B", x"F052", x"EC76", x"EAEA", x"EB13", x"EC5A", x"EDD4", x"EF48",
		x"F0B6", x"F227", x"F3B1", x"F554", x"F747", x"F995", x"FC1E", x"FEC7",
		x"016D", x"0424", x"06E4", x"09B6", x"0C62", x"0EA2", x"1077", x"11E6",
		x"1312", x"13EE", x"148C", x"14D7", x"14F1", x"1505", x"14DC", x"1478",
		x"13BC", x"127F", x"1029", x"0C85", x"07B2", x"01C8", x"FB91", x"F59F",
		x"F088", x"ED26", x"EC35", x"EE80", x"F415", x"FC56", x"057B", x"0D82",
		x"12D1", x"1493", x"13A4", x"118A", x"0FE7", x"0FC4", x"1126", x"12E0",
		x"1346", x"10E4", x"0B73", x"0414", x"FC71", x"F5F6", x"F159", x"EE96",
		x"ED3E", x"ECF6", x"ECBB", x"EC56", x"EBB7", x"EBBB", x"ED7C", x"F21D",
		x"F97B", x"022A", x"0A4C", x"1079", x"141D", x"15C4", x"1580", x"1339",
		x"0EC4", x"085B", x"0088", x"F88A", x"F1A5", x"ECEC", x"EAA2", x"EA50",
		x"EAA1", x"EB17", x"EB75", x"EC4B", x"EE48", x"F1C1", x"F70F", x"FE01",
		x"05B9", x"0CC4", x"11B6", x"1394", x"12A3", x"1042", x"0E33", x"0DF4",
		x"0F9C", x"1212", x"137D", x"1251", x"0DF6", x"0726", x"FF66", x"F858",
		x"F2CC", x"EF3E", x"ED1D", x"EBFE", x"EB82", x"EB3D", x"EB3D", x"EB55",
		x"EBBE", x"EC94", x"EDE9", x"EFDF", x"F253", x"F489", x"F5E1", x"F588",
		x"F37B", x"F076", x"ED79", x"EC1C", x"ED96", x"F238", x"F924", x"00CC",
		x"07B3", x"0D18", x"1107", x"1389", x"14F1", x"1596", x"15BD", x"1593",
		x"14C8", x"1290", x"0E70", x"084A", x"0088", x"F886", x"F1A3", x"ECD8",
		x"EA7A", x"EA1B", x"EA8B", x"EB2F", x"EBE2", x"ECE9", x"EE7F", x"F061",
		x"F1DB", x"F274", x"F1E6", x"F035", x"EE2B", x"EC66", x"EB88", x"EB5F",
		x"EB4F", x"EB41", x"EBB1", x"EDA5", x"F1D9", x"F864", x"005E", x"0882",
		x"0F00", x"1312", x"14CA", x"14F1", x"145D", x"13A6", x"12F6", x"123B",
		x"114A", x"0FEF", x"0E1D", x"0BFC", x"09B6", x"075B", x"04DC", x"023D",
		x"FF6C", x"FCA6", x"F9D7", x"F744", x"F4BC", x"F211", x"EF93", x"ED7A",
		x"EC07", x"EB51", x"EB3A", x"EBA0", x"EC97", x"EE3A", x"F060", x"F2D7",
		x"F53A", x"F6E2", x"F738", x"F5EB", x"F31D", x"EFD5", x"ED28", x"EC59",
		x"EE37", x"F333", x"FADF", x"03D1", x"0C19", x"11B9", x"139D", x"11C2",
		x"0D32", x"0794", x"0285", x"FF71", x"FF6B", x"0265", x"07BB", x"0D5C",
		x"1199", x"12E6", x"10BF", x"0BF9", x"05DD", x"0019", x"FB9C", x"F8B7",
		x"F72C", x"F68A", x"F5E5", x"F49E", x"F283", x"F01B", x"EDE2", x"EC40",
		x"EB42", x"EAFA", x"EB25", x"EB25", x"EAE7", x"EAD0", x"EC05", x"EF9A",
		x"F595", x"FD40", x"0547", x"0C2C", x"10FC", x"139A", x"14A2", x"14D4",
		x"149C", x"13C6", x"11FA", x"0EFA", x"0A89", x"0498", x"FD8B", x"F63A",
		x"F054", x"ED2D", x"ED7C", x"F037", x"F3E9", x"F660", x"F669", x"F3EB",
		x"F04A", x"ED67", x"ED83", x"F147", x"F792", x"FE2C", x"02F5", x"04DA",
		x"0409", x"010D", x"FD09", x"F8CD", x"F4EC", x"F22A", x"F0B0", x"F062",
		x"F0DE", x"F205", x"F3E4", x"F68C", x"FA0C", x"FE3C", x"032F", x"089F",
		x"0DE4", x"122D", x"1427", x"1354", x"0F99", x"09F1", x"0359", x"FD28",
		x"F7EE", x"F3CD", x"F0DB", x"EED9", x"EDB4", x"ED53", x"ED35", x"ED4A",
		x"ED91", x"EE50", x"EFDF", x"F24C", x"F54F", x"F856", x"FAAD", x"FBF8",
		x"FBC0", x"F9F7", x"F6FE", x"F363", x"F02D", x"EDDC", x"EC8F", x"EC5D",
		x"EDC0", x"F17A", x"F7BE", x"FFC2", x"07FD", x"0EB9", x"131E", x"1559",
		x"15E6", x"159A", x"146D", x"1207", x"0DA4", x"06F9", x"FE7D", x"F60F",
		x"EFA5", x"EBE1", x"EA9E", x"EAB9", x"EB9E", x"ECB2", x"ED9A", x"EE2C",
		x"EE43", x"EDF5", x"ED72", x"ECBE", x"EC07", x"EB61", x"EB02", x"EB0B",
		x"EB88", x"EC98", x"EE3C", x"F09F", x"F34C", x"F613", x"F880", x"FA90",
		x"FBCD", x"FC26", x"FB9F", x"F9FD", x"F777", x"F467", x"F188", x"EF0F",
		x"ED80", x"ECFD", x"EE36", x"F1C0", x"F7D2", x"FF9F", x"077A", x"0E44",
		x"12AA", x"149F", x"14C7", x"1446", x"1402", x"1445", x"149E", x"147E",
		x"13CC", x"132B", x"134B", x"13F4", x"1496", x"13CB", x"109B", x"0ACA",
		x"02FA", x"FAC9", x"F3BA", x"EEEC", x"EC34", x"EB03", x"EABC", x"EAD7",
		x"EB1B", x"EB52", x"EBB3", x"ECB7", x"EE49", x"F06E", x"F2D2", x"F582",
		x"F84E", x"FAF9", x"FD02", x"FE0C", x"FDF4", x"FCC5", x"FAC5", x"F838",
		x"F56A", x"F29B", x"F024", x"EE2A", x"ECE0", x"EC4D", x"EBD2", x"EB7C",
		x"EB22", x"EAFA", x"EB54", x"ECA5", x"EF0F", x"F2B3", x"F7D2", x"FDF4",
		x"04CB", x"0B58", x"10A1", x"1386", x"1323", x"0F46", x"0872", x"0033",
		x"F7FF", x"F16C", x"ED56", x"EB82", x"EB35", x"EBAC", x"EC37", x"EC97",
		x"EC90", x"EC1C", x"EB68", x"EB3E", x"EC4E", x"EF06", x"F348", x"F8E9",
		x"FF8A", x"065A", x"0C92", x"115A", x"13B9", x"1306", x"0EB3", x"072B",
		x"FE10", x"F57C", x"EF33", x"EBF1", x"EB17", x"EB38", x"EB69", x"EB93",
		x"EC72", x"EF1F", x"F447", x"FBC8", x"041F", x"0B68", x"1001", x"11A4",
		x"10E6", x"0EA1", x"0BA1", x"07EF", x"0483", x"0226", x"0189", x"0353",
		x"072C", x"0C23", x"10B7", x"136F", x"131E", x"0F4F", x"088A", x"0022",
		x"F7CB", x"F120", x"ED2D", x"EC74", x"EE87", x"F26F", x"F6D4", x"FA73",
		x"FC85", x"FCD4", x"FBA2", x"F963", x"F66A", x"F329", x"F030", x"EDE7",
		x"EC56", x"EB53", x"EAF9", x"EB3D", x"EBCE", x"EC70", x"ECDB", x"ED24",
		x"ED76", x"EDAF", x"ED9F", x"ED11", x"EC5B", x"EBB1", x"EB51", x"EBB2",
		x"ED61", x"F13B", x"F774", x"FF5A", x"075C", x"0E17", x"1299", x"14C0",
		x"1530", x"14EF", x"14CA", x"14F0", x"14DC", x"1436", x"130F", x"120F",
		x"11E7", x"12BC", x"13F4", x"140B", x"11F6", x"0CC6", x"0554", x"FD67",
		x"F6A8", x"F227", x"EFE4", x"EF28", x"EF8A", x"F0E8", x"F350", x"F6DA",
		x"FB8E", x"013C", x"078B", x"0D8F", x"1205", x"13D0", x"1284", x"0E88",
		x"0924", x"03AA", x"FF79", x"FD53", x"FD3A", x"FF33", x"026B", x"065C",
		x"0A2D", x"0D6D", x"100D", x"1203", x"138A", x"148F", x"1519", x"154A",
		x"154A", x"1535", x"14C4", x"1406", x"12C2", x"1152", x"0FE8", x"0EC0",
		x"0D63", x"0B09", x"0782", x"0275", x"FC53", x"F5DC", x"F04C", x"ECFF",
		x"ECC5", x"EFB0", x"F47B", x"F9D3", x"FEAC", x"020B", x"0410", x"0536",
		x"062B", x"07C6", x"0A60", x"0DC8", x"10F2", x"12D1", x"1227", x"0E7B",
		x"0869", x"015E", x"FAAC", x"F5FE", x"F450", x"F5E9", x"FA30", x"0056",
		x"074F", x"0DB6", x"120F", x"12A9", x"0F0E", x"07B6", x"FE8D", x"F5D8",
		x"EF6A", x"EC0D", x"EB55", x"EC3D", x"ED3D", x"ED88", x"ECE6", x"EC28",
		x"ECA9", x"EFF8", x"F613", x"FE62", x"071F", x"0E67", x"12E1", x"13CE",
		x"118C", x"0CD7", x"06D0", x"007C", x"FA7C", x"F514", x"F0A4", x"ED6C",
		x"EB9C", x"EB0B", x"EB2B", x"EB60", x"EB4E", x"EAF5", x"EB19", x"ECC7",
		x"F07E", x"F635", x"FD74", x"053D", x"0C5C", x"11CF", x"1503", x"15EC",
		x"1580", x"14A8", x"13E5", x"1332", x"124A", x"10A2", x"0DC7", x"0997",
		x"03E6", x"FD2B", x"F63D", x"F0A6", x"ED52", x"ED04", x"F01D", x"F60D",
		x"FE0D", x"0667", x"0D9E", x"1255", x"1465", x"1446", x"129B", x"109D",
		x"0F14", x"0E94", x"0F34", x"10A5", x"1251", x"13BB", x"1474", x"13F4",
		x"11CF", x"0DFF", x"0866", x"0178", x"F9EE", x"F313", x"EE54", x"EC6B",
		x"ED9D", x"F166", x"F728", x"FDE4", x"0505", x"0B8E", x"10CA", x"13D9",
		x"13C7", x"105E", x"09BC", x"0146", x"F8C3", x"F1C8", x"ED36", x"EADD",
		x"EA0B", x"EA3D", x"EB0A", x"EC18", x"ED43", x"EE8E", x"EFD1", x"F0B5",
		x"F0D2", x"EFDE", x"EE1C", x"EC80", x"EC3E", x"EE96", x"F406", x"FBEE",
		x"04AA", x"0C76", x"11A4", x"1310", x"1091", x"0B39", x"04A3", x"FE62",
		x"F9C8", x"F7AA", x"F8A8", x"FCC5", x"0301", x"09F7", x"0FC0", x"1302",
		x"12F9", x"0FF7", x"0B0D", x"05BD", x"011B", x"FDC9", x"FBD2", x"FAC9",
		x"FA3B", x"F9EF", x"F9AF", x"F9D8", x"FA47", x"FB34", x"FCD1", x"FF2B",
		x"0289", x"06DF", x"0BEE", x"107B", x"136D", x"136D", x"107A", x"0B32",
		x"04F3", x"FED8", x"F9D7", x"F672", x"F4CB", x"F4C2", x"F60D", x"F849",
		x"FB82", x"FFDD", x"054C", x"0B35", x"1049", x"134A", x"1322", x"0FC6",
		x"09F6", x"0363", x"FD78", x"F993", x"F818", x"F8D5", x"FB81", x"FF72",
		x"03A4", x"074E", x"09A7", x"0A11", x"07F3", x"02F4", x"FBFA", x"F4AF",
		x"EF4D", x"ECE7", x"ED93", x"F016", x"F2E4", x"F4D1", x"F527", x"F420",
		x"F215", x"EFC2", x"ED9E", x"EBFB", x"EB94", x"ECEF", x"F09C", x"F677",
		x"FDA3", x"0536", x"0BFA", x"1120", x"141D", x"1524", x"1479", x"12F4",
		x"1133", x"0FC1", x"0EB0", x"0DB7", x"0C92", x"0B10", x"08D8", x"0613",
		x"02FD", x"0010", x"FD56", x"FAD4", x"F871", x"F62C", x"F447", x"F292",
		x"F11D", x"EFA5", x"EE61", x"ED13", x"EBD3", x"EB1E", x"EB79", x"ED89",
		x"F1A7", x"F7D5", x"FF7D", x"0756", x"0E16", x"1283", x"13DD", x"123F",
		x"0E3E", x"0889", x"01CE", x"FAC5", x"F45B", x"EF47", x"EC7D", x"ED1C",
		x"F181", x"F900", x"01C9", x"09CA", x"0FBA", x"1351", x"14D6", x"1497",
		x"12C3", x"0F4B", x"09F4", x"030F", x"FB39", x"F3F3", x"EEF7", x"EDAD",
		x"F0B3", x"F768", x"0015", x"0893", x"0F3E", x"1389", x"158F", x"15FD",
		x"14D5", x"11A0", x"0C34", x"0515", x"FD29", x"F59A", x"EF81", x"EBD2",
		x"EAEE", x"ECAC", x"F0BB", x"F709", x"FF14", x"07C4", x"0F2D", x"13C7",
		x"1530", x"1465", x"12D5", x"117C", x"10B4", x"100B", x"0EE5", x"0C90",
		x"086B", x"0281", x"FB6F", x"F496", x"EF48", x"ECB2", x"ED08", x"EFE9",
		x"F453", x"F8FC", x"FD4E", x"00D3", x"03C7", x"0648", x"088B", x"0A9C",
		x"0C47", x"0DA9", x"0ED9", x"0FF3", x"1120", x"1245", x"1371", x"145A",
		x"14D8", x"1437", x"119B", x"0C4A", x"04DE", x"FC64", x"F4BB", x"EEFD",
		x"EBA9", x"EA33", x"EA11", x"EB08", x"ED46", x"F1A5", x"F88D", x"0145",
		x"09EA", x"1098", x"13CB", x"132E", x"0F8A", x"09FE", x"0370", x"FCB4",
		x"F64C", x"F0BD", x"ED1E", x"ECC7", x"F039", x"F6F9", x"FF72", x"0791",
		x"0E07", x"1230", x"13F6", x"1339", x"1009", x"0A31", x"02AC", x"FA9E",
		x"F35C", x"EE2D", x"EB5E", x"EA80", x"EAB1", x"EAFC", x"EB23", x"EB9E",
		x"ECEE", x"EEB2", x"F006", x"F013", x"EEE2", x"ED33", x"EC4A", x"EDC1",
		x"F23E", x"F987", x"021D", x"0A30", x"1030", x"1343", x"132C", x"104F",
		x"0B04", x"0456", x"FD6A", x"F753", x"F281", x"EF2E", x"ED19", x"EBED",
		x"EB67", x"EB1E", x"EAE5", x"EADD", x"EB20", x"EBE4", x"ED53", x"EF83",
		x"F229", x"F488", x"F67D", x"F7C7", x"F888", x"F8A8", x"F834", x"F709",
		x"F5C0", x"F430", x"F237", x"EFA6", x"ED18", x"EB9C", x"EC77", x"F05A",
		x"F6D7", x"FEB5", x"06AE", x"0D86", x"1237", x"13E8", x"1217", x"0CED",
		x"054D", x"FCF4", x"F565", x"EF7F", x"EBC0", x"E9ED", x"E9DE", x"EB47",
		x"EE48", x"F334", x"FA23", x"029B", x"0AA6", x"10CE", x"1433", x"1556",
		x"151E", x"1444", x"12F7", x"10F2", x"0DD0", x"0965", x"03D8", x"FD83",
		x"F701", x"F162", x"EDB3", x"ECCA", x"EEEA", x"F2EE", x"F6E4", x"F97B",
		x"F9FF", x"F8E0", x"F691", x"F3B1", x"F0E9", x"EE97", x"ED0D", x"EC6F",
		x"EC8F", x"ED1F", x"EE5E", x"F00C", x"F240", x"F4E1", x"F7F2", x"FB7E",
		x"FF46", x"0347", x"072A", x"0A95", x"0D33", x"0EDB", x"0F9A", x"0F29",
		x"0D05", x"08B2", x"024F", x"FAC6", x"F3DB", x"EEAC", x"EC48", x"ECBF",
		x"EF6A", x"F2FC", x"F654", x"F8C9", x"FA9E", x"FBF0", x"FD6D", x"FF4B",
		x"01DD", x"0523", x"08C4", x"0C82", x"0FC0", x"1213", x"1353", x"13B1",
		x"12E6", x"10E4", x"0D3B", x"0788", x"008B", x"F914", x"F25A", x"ED99",
		x"EBB6", x"EC85", x"EF6C", x"F344", x"F70A", x"FA4C", x"FC88", x"FD6A",
		x"FCCF", x"FAAE", x"F75E", x"F352", x"EF60", x"ECC0", x"EC8B", x"EF45",
		x"F4EF", x"FCD7", x"058A", x"0D22", x"1219", x"138E", x"11D3", x"0DC4",
		x"08CA", x"046B", x"01B8", x"013D", x"02A2", x"053B", x"085F", x"0B91",
		x"0E4A", x"0FEC", x"0FDF", x"0D97", x"08CB", x"01F9", x"FA1F", x"F2F6",
		x"EDF7", x"EC13", x"ECFC", x"EF70", x"F20E", x"F420", x"F579", x"F668",
		x"F7BE", x"FA00", x"FDEA", x"033F", x"0973", x"0EFF", x"12A3", x"1347",
		x"10C9", x"0C22", x"06DB", x"02E1", x"0109", x"0154", x"0334", x"05FD",
		x"092E", x"0C31", x"0EAC", x"106A", x"1165", x"1175", x"10D2", x"0F5F",
		x"0D4D", x"0A43", x"0671", x"01A0", x"FC3F", x"F6B1", x"F18F", x"EDAE",
		x"EBE5", x"ECD3", x"F07C", x"F692", x"FE53", x"0654", x"0D83", x"126F",
		x"145B", x"132D", x"0FAD", x"0A98", x"0513", x"FFBB", x"FAE4", x"F728",
		x"F487", x"F2D3", x"F1AE", x"F086", x"EF2B", x"EDB3", x"EC48", x"EB80",
		x"EB74", x"EC0C", x"ECDB", x"ED4C", x"ED2C", x"EC8C", x"EC1B", x"ED00",
		x"F051", x"F630", x"FDD1", x"05BD", x"0C49", x"1022", x"1038", x"0C1A",
		x"04C2", x"FC0F", x"F481", x"EF64", x"EC70", x"EAFD", x"EA5B", x"EAA9",
		x"EC63", x"F031", x"F65D", x"FE72", x"06EE", x"0DE2", x"118E", x"10EB",
		x"0C63", x"051C", x"FCA0", x"F4C0", x"EED6", x"EB8D", x"EAE1", x"EBC6",
		x"ECB0", x"ECCC", x"EC39", x"EBAC", x"EBD6", x"EC8F", x"ED48", x"ED91",
		x"ED54", x"ECBA", x"EBDB", x"EB3D", x"EB05", x"EB10", x"EB65", x"EBB0",
		x"EBC4", x"EB85", x"EB2C", x"EAE6", x"EAE1", x"EB66", x"EC6F", x"EDBA",
		x"EF61", x"F15C", x"F353", x"F56A", x"F793", x"F9DE", x"FC79", x"FF7C",
		x"029D", x"05DA", x"0919", x"0C1C", x"0EC9", x"10C9", x"1213", x"12A8",
		x"12D2", x"123E", x"10FB", x"0F4B", x"0D52", x"0B2C", x"08D4", x"06A3",
		x"04B6", x"03A1", x"03C1", x"04E9", x"06D5", x"094A", x"0C36", x"0F48",
		x"11F0", x"13B6", x"1418", x"12A8", x"0F32", x"09AD", x"0290", x"FABB",
		x"F38C", x"EE77", x"EC57", x"ED8B", x"F1DD", x"F85F", x"FFBC", x"06DA",
		x"0CA8", x"10D2", x"1377", x"14C1", x"1505", x"14CC", x"1433", x"1390",
		x"12BC", x"11B1", x"1071", x"0F3B", x"0DF4", x"0C8E", x"0AFC", x"08C2",
		x"05BB", x"0188", x"FC22", x"F63F", x"F0D3", x"ED67", x"ED2D", x"F073",
		x"F601", x"FB97", x"FF1C", x"FF23", x"FB6B", x"F564", x"EFD4", x"ED35",
		x"EE8B", x"F2BB", x"F6B3", x"F836", x"F668", x"F276", x"EED0", x"EE0C",
		x"F13F", x"F739", x"FD5F", x"009C", x"FF6D", x"FA76", x"F3E6", x"EED1",
		x"ED25", x"EF28", x"F2E2", x"F5E6", x"F688", x"F433", x"F073", x"ED80",
		x"ED86", x"F11B", x"F73A", x"FDC9", x"02B1", x"04C7", x"03EE", x"00C8",
		x"FCB6", x"F885", x"F50A", x"F296", x"F147", x"F131", x"F213", x"F3F9",
		x"F6AA", x"F9E3", x"FD53", x"00C4", x"0405", x"06F2", x"096B", x"0B8C",
		x"0D67", x"0F39", x"10F5", x"1279", x"13C5", x"14BA", x"1559", x"1573",
		x"1520", x"14A7", x"13D5", x"12C6", x"1146", x"0F63", x"0D02", x"0A2A",
		x"06F6", x"039E", x"0063", x"FDBE", x"FBF4", x"FB5D", x"FBFA", x"FDE9",
		x"00D7", x"044E", x"0798", x"0A61", x"0C61", x"0D46", x"0C3B", x"08C7",
		x"0329", x"FC39", x"F55B", x"EFEC", x"ED34", x"EDD9", x"F1BB", x"F818",
		x"FF85", x"06EC", x"0D1A", x"1174", x"1362", x"12D1", x"0FB0", x"0A4B",
		x"0340", x"FB62", x"F421", x"EEB0", x"EBF2", x"EBFE", x"EE1B", x"F15A",
		x"F4F1", x"F82C", x"FB18", x"FD5B", x"FF5C", x"012C", x"032F", x"0593",
		x"0865", x"0BAE", x"0EEE", x"11BD", x"138D", x"148A", x"14FB", x"14B0",
		x"1304", x"0F03", x"0867", x"0026", x"F7E9", x"F156", x"ECDE", x"EA6F",
		x"E9A4", x"EA1F", x"EC17", x"EFB2", x"F58E", x"FD5D", x"061D", x"0DD3",
		x"1258", x"12A2", x"0E8F", x"0733", x"FEA5", x"F6D8", x"F11E", x"ED86",
		x"EBF4", x"EC5B", x"EEF5", x"F3DE", x"FABD", x"02B0", x"0A67", x"1084",
		x"141A", x"156D", x"156A", x"1515", x"148C", x"13A8", x"121C", x"1030",
		x"0E5E", x"0D8B", x"0E10", x"0F9C", x"11C4", x"13AB", x"14E0", x"155D",
		x"157B", x"154F", x"149D", x"12C0", x"0F20", x"096B", x"0200", x"FA1C",
		x"F301", x"EE22", x"EB77", x"EAFD", x"EBA4", x"ECDA", x"EE1E", x"EF2A",
		x"EFF7", x"F10E", x"F296", x"F4A9", x"F771", x"FAE9", x"FED8", x"02A6",
		x"059A", x"0784", x"0860", x"0800", x"063E", x"0344", x"FF7F", x"FBB4",
		x"F878", x"F62F", x"F514", x"F55C", x"F721", x"F9E0", x"FD40", x"00B9",
		x"03DB", x"0643", x"0763", x"069C", x"03AD", x"FEB4", x"F8B3", x"F2B8",
		x"EE3A", x"EC64", x"EDF0", x"F30E", x"FACC", x"0379", x"0B6F", x"113F",
		x"143E", x"1455", x"1244", x"0F58", x"0CC6", x"0B2F", x"0B15", x"0C2F",
		x"0E13", x"1034", x"1228", x"13B3", x"1486", x"1490", x"13E4", x"12FC",
		x"122D", x"117E", x"10AA", x"0F44", x"0D1F", x"0A0B", x"0630", x"01E7",
		x"FDAE", x"F9F2", x"F718", x"F581", x"F5B3", x"F845", x"FD29", x"03CB",
		x"0AE8", x"10B1", x"1388", x"1323", x"1092", x"0D9A", x"0BBC", x"0BD0",
		x"0DB0", x"1042", x"12A1", x"142E", x"152C", x"15C1", x"1530", x"127E",
		x"0CB8", x"04B2", x"FC01", x"F44F", x"EEC2", x"EB9D", x"EADE", x"EC14",
		x"EF47", x"F486", x"FBB5", x"0401", x"0BE3", x"11A6", x"1480", x"1494",
		x"12FC", x"10FB", x"0F33", x"0DDE", x"0CB6", x"0BD4", x"0B3B", x"0B4F",
		x"0C07", x"0D16", x"0EB2", x"1074", x"1226", x"1381", x"1492", x"150D",
		x"1507", x"148D", x"13DB", x"135B", x"12C3", x"1199", x"0FA3", x"0CFF",
		x"09D9", x"0641", x"026D", x"FE6E", x"FAF5", x"F86B", x"F75F", x"F82E",
		x"FB53", x"00EC", x"07D2", x"0E2C", x"120E", x"12B2", x"10A4", x"0D9B",
		x"0B2D", x"0A3D", x"0B24", x"0D3F", x"0FEE", x"1252", x"13FD", x"14B9",
		x"1490", x"133D", x"1069", x"0BB1", x"054E", x"FD8C", x"F5A0", x"EF55",
		x"EC2E", x"ECDA", x"F10B", x"F7C7", x"FF9D", x"071B", x"0D5E", x"11B4",
		x"13EF", x"1468", x"137A", x"11B4", x"0F8B", x"0D70", x"0BC2", x"0A9E",
		x"09FD", x"09D8", x"0A1B", x"0AD3", x"0C42", x"0E42", x"1053", x"1249",
		x"13B3", x"148E", x"14EF", x"14F1", x"14AB", x"146E", x"1436", x"13A5",
		x"124A", x"0F9C", x"0B20", x"04B0", x"FCBE", x"F4D8", x"EED9", x"EBF9",
		x"EC18", x"ED8F", x"EEAD", x"EE7F", x"ED7C", x"ECF9", x"EEBA", x"F3DF",
		x"FB79", x"03B8", x"0A28", x"0D58", x"0D68", x"0B3C", x"0785", x"0334",
		x"FEF4", x"FBE4", x"FAC8", x"FC13", x"FFD1", x"0540", x"0B5A", x"1070",
		x"1315", x"1264", x"0E61", x"07BF", x"FF83", x"F741", x"F091", x"ECAE",
		x"EC05", x"EE14", x"F1AF", x"F534", x"F76B", x"F7B7", x"F66B", x"F407",
		x"F130", x"EEA8", x"ECD2", x"EBB7", x"EB5C", x"EBA7", x"EC8F", x"EE12",
		x"F043", x"F2B6", x"F533", x"F746", x"F86F", x"F88D", x"F7F6", x"F6C5",
		x"F519", x"F2FD", x"F094", x"EE0F", x"EC1D", x"EB8D", x"ED23", x"F155",
		x"F7E8", x"FFB5", x"0750", x"0D82", x"11A3", x"13C4", x"1439", x"138F",
		x"11F0", x"0F9D", x"0CDE", x"0A07", x"07C2", x"067E", x"06A0", x"07E8",
		x"0A22", x"0CCB", x"0F4A", x"1153", x"129C", x"133A", x"1384", x"1399",
		x"1382", x"1304", x"11DE", x"0FCD", x"0C93", x"07E5", x"01E6", x"FAF7",
		x"F43C", x"EF07", x"EC87", x"ECF6", x"EFA3", x"F37B", x"F71A", x"F994",
		x"FA7D", x"F9CA", x"F7A2", x"F4B6", x"F1C6", x"EEE7", x"EC99", x"EB13",
		x"EA57", x"EA54", x"EAE1", x"EBAC", x"ECA2", x"ED98", x"EE56", x"EEAF",
		x"EEA7", x"EE67", x"EDDE", x"ED22", x"EC42", x"EB73", x"EB90", x"ED26",
		x"F0E2", x"F6EF", x"FE88", x"0673", x"0D1D", x"11CA", x"1419", x"14B5",
		x"1487", x"142B", x"13F2", x"140C", x"1486", x"14DC", x"147A", x"1256",
		x"0E11", x"07A3", x"0005", x"F853", x"F1E2", x"ED92", x"EBB9", x"EBDB",
		x"ED22", x"EE80", x"EF57", x"EF3C", x"EE28", x"ECA0", x"EBA2", x"EC25",
		x"EE4F", x"F0D6", x"F209", x"F101", x"EEBA", x"ED39", x"EE11", x"F123",
		x"F555", x"F946", x"FBEB", x"FCDE", x"FC1D", x"F9FB", x"F6C8", x"F2F2",
		x"EF5E", x"ECAF", x"EBA3", x"ECC0", x"F058", x"F624", x"FD4C", x"04CA",
		x"0B5D", x"1055", x"1345", x"14A9", x"14E1", x"14CA", x"1485", x"1442",
		x"13C8", x"1285", x"0FCD", x"0B2C", x"04BC", x"FD05", x"F585", x"EF99",
		x"EC55", x"EBD6", x"ED68", x"EFF8", x"F288", x"F4A2", x"F651", x"F7D5",
		x"F9AA", x"FC58", x"0020", x"04F2", x"0A6A", x"0F9A", x"132D", x"1412",
		x"11EF", x"0D01", x"05FB", x"FDF1", x"F625", x"EFEC", x"EC32", x"EB4A",
		x"ED1D", x"F150", x"F763", x"FE97", x"05FF", x"0C99", x"1155", x"1387",
		x"1301", x"0FCF", x"0A81", x"0396", x"FC04", x"F4F2", x"EF68", x"EC65",
		x"EC26", x"EEA5", x"F38F", x"FA26", x"0190", x"088D", x"0E57", x"125C",
		x"141E", x"134F", x"0FBF", x"0988", x"01AE", x"F96D", x"F246", x"ED9B",
		x"EC87", x"EEDD", x"F322", x"F791", x"FA6E", x"FAA7", x"F81D", x"F3C9",
		x"EF6D", x"ECDD", x"ED82", x"F1A9", x"F88F", x"00C7", x"08D2", x"0F46",
		x"134F", x"1446", x"1278", x"0E2B", x"080F", x"00FA", x"F9DB", x"F361",
		x"EE9B", x"EC60", x"ECC4", x"EFE1", x"F55C", x"FC7C", x"0424", x"0B31",
		x"10AC", x"13DF", x"1461", x"1223", x"0D3B", x"0645", x"FE1F", x"F629",
		x"F009", x"ECFC", x"EDB6", x"F17C", x"F68B", x"FAC1", x"FC4F", x"FA87",
		x"F615", x"F0F9", x"ED8B", x"ED67", x"F06C", x"F4EA", x"F8AA", x"F9E0",
		x"F806", x"F3FB", x"EFA8", x"ED17", x"EE05", x"F2AE", x"FA23", x"02A2",
		x"0A8D", x"1062", x"13B3", x"144E", x"1230", x"0DC7", x"076D", x"FFF0",
		x"F841", x"F1B1", x"ED76", x"EC24", x"EDE4", x"F1C8", x"F6F4", x"FC79",
		x"0198", x"0628", x"09D5", x"0CB4", x"0EC4", x"1063", x"117D", x"126A",
		x"133E", x"13C9", x"1431", x"1478", x"14BE", x"14B4", x"142F", x"12D8",
		x"1045", x"0C1D", x"068B", x"FFCD", x"F8B3", x"F24C", x"EDE2", x"EC48",
		x"EE07", x"F2A0", x"F957", x"00B9", x"07F5", x"0E08", x"1226", x"13DF",
		x"12E5", x"0EEE", x"0813", x"FF69", x"F6CA", x"F041", x"ECB3", x"EBB3",
		x"EBD5", x"EC10", x"EC26", x"EC7F", x"EE4F", x"F28A", x"F968", x"01C5",
		x"098F", x"0E30", x"0E49", x"09D6", x"0230", x"F9C8", x"F2BA", x"EE29",
		x"EC41", x"EBD7", x"EBFC", x"EC2B", x"ECF1", x"EF22", x"F3B3", x"FACE",
		x"02EC", x"0A1A", x"0DF6", x"0D7A", x"091D", x"023F", x"FA77", x"F367",
		x"EE76", x"EC80", x"ED98", x"F0DC", x"F4D4", x"F834", x"FA98", x"FC35",
		x"FDB6", x"FF4E", x"0127", x"0347", x"05DD", x"08A2", x"0B78", x"0DE8",
		x"0FE5", x"117B", x"12BD", x"13B3", x"1461", x"1497", x"148B", x"1450",
		x"13C8", x"12D1", x"115F", x"0FA7", x"0DF4", x"0C72", x"0B22", x"0A12",
		x"08EC", x"071A", x"03CB", x"FF22", x"F96E", x"F3C3", x"EF51", x"ED8F",
		x"EF22", x"F3A5", x"F97E", x"FE5D", x"006B", x"FEBF", x"F9EA", x"F3B9",
		x"EEC1", x"ECF4", x"EE89", x"F226", x"F585", x"F6D4", x"F56B", x"F1E6",
		x"EE57", x"ED15", x"EF88", x"F59B", x"FDE2", x"066A", x"0D97", x"1275",
		x"1477", x"13F8", x"10F9", x"0BCB", x"04D2", x"FCDD", x"F557", x"EFAD",
		x"ECF3", x"ED97", x"F122", x"F68F", x"FC3A", x"00B1", x"0310", x"0356",
		x"01FB", x"FFA0", x"FCE7", x"F9EF", x"F712", x"F48F", x"F2C4", x"F211",
		x"F272", x"F3D8", x"F643", x"F992", x"FD99", x"0226", x"0720", x"0C18",
		x"1058", x"131A", x"13CB", x"122A", x"0DEA", x"073B", x"FF12", x"F6F0",
		x"F07D", x"ECDB", x"EC97", x"EF0C", x"F38E", x"F956", x"FF5C", x"04F5",
		x"09A4", x"0D3D", x"0FD6", x"11A7", x"12F9", x"13DB", x"1463", x"144C",
		x"13B3", x"12A2", x"1113", x"0EAB", x"0B97", x"08D8", x"0768", x"0819",
		x"0AC2", x"0E7F", x"11C2", x"12AC", x"1002", x"0A23", x"0311", x"FDBA",
		x"FC29", x"FF07", x"0524", x"0C0C", x"111A", x"129A", x"10F3", x"0DE5",
		x"0BDE", x"0C18", x"0E6E", x"1128", x"121C", x"0FB2", x"0A14", x"0331",
		x"FD26", x"F994", x"F8D2", x"FA81", x"FDB6", x"01E9", x"060B", x"097B",
		x"0B9E", x"0C34", x"0B71", x"0980", x"06A4", x"030F", x"FF59", x"FC3E",
		x"FA2F", x"F960", x"F9CD", x"FB92", x"FE2B", x"01A1", x"04F0", x"07C0",
		x"09BB", x"0ABF", x"0B08", x"0A79", x"0923", x"0706", x"0437", x"00DE",
		x"FD55", x"FA01", x"F6CA", x"F3E5", x"F141", x"EEF8", x"ED6A", x"EC57",
		x"EBBC", x"EB47", x"EB02", x"EAEE", x"EB3E", x"EC21", x"ED8D", x"EF86",
		x"F1CF", x"F3FA", x"F57E", x"F621", x"F5C8", x"F459", x"F23D", x"EFFA",
		x"EDC4", x"EC22", x"EAF5", x"EA77", x"EA9C", x"EAFB", x"EB70", x"EBDA",
		x"EC9E", x"EE25", x"F0EF", x"F4F5", x"FA86", x"0115", x"07F4", x"0E08",
		x"1219", x"13A8", x"1291", x"0F81", x"0B72", x"071E", x"030B", x"FFB7",
		x"FCDC", x"FA8E", x"F88F", x"F6E3", x"F582", x"F45C", x"F328", x"F1D5",
		x"F035", x"EE5A", x"ECBE", x"EBA1", x"EB77", x"EC76", x"EEF0", x"F30D",
		x"F8E3", x"0004", x"079C", x"0E51", x"129C", x"1337", x"0F6C", x"0844",
		x"FF9A", x"F790", x"F16B", x"EDA9", x"EBBE", x"EB52", x"EC31", x"EE86",
		x"F2BE", x"F918", x"0114", x"0956", x"0FB8", x"12B2", x"1156", x"0BD2",
		x"038F", x"FAEF", x"F3B3", x"EEBC", x"EBDB", x"EAA5", x"EB4B", x"EDFF",
		x"F310", x"FA31", x"026D", x"0A64", x"10B2", x"1473", x"158D", x"143A",
		x"10CC", x"0B5F", x"0410", x"FBAF", x"F3E0", x"EE1D", x"EB42", x"EA8A",
		x"EAA2", x"EACB", x"EB0D", x"EBE0", x"ED82", x"F065", x"F49F", x"FA2B",
		x"00F6", x"081F", x"0E76", x"1261", x"135A", x"119E", x"0DEC", x"0989",
		x"0532", x"015F", x"FE4A", x"FBD3", x"F9C7", x"F806", x"F660", x"F479",
		x"F2A9", x"F0E9", x"EF84", x"EE41", x"ECF7", x"EBD9", x"EAFE", x"EAB6",
		x"EB0A", x"EBEB", x"ED4E", x"EF5C", x"F1C5", x"F3E7", x"F52F", x"F51F",
		x"F3D1", x"F140", x"EE44", x"EC5A", x"ECCD", x"F04C", x"F6C7", x"FEE4",
		x"071D", x"0DF9", x"1285", x"1462", x"13AA", x"10C3", x"0BA7", x"04B8",
		x"FCB0", x"F4D7", x"EF28", x"ECD5", x"EEA9", x"F38F", x"F9D6", x"FFAE",
		x"0363", x"0401", x"0162", x"FC44", x"F5FB", x"F05B", x"ECFD", x"EC9C",
		x"EF5C", x"F45B", x"FA83", x"00A4", x"05F7", x"09E4", x"0C47", x"0D70",
		x"0D3F", x"0B44", x"073E", x"013A", x"FA08", x"F31C", x"EE31", x"EC0D",
		x"EC97", x"EE32", x"EF52", x"EF0B", x"EDC7", x"ECF1", x"EEB6", x"F3AA",
		x"FB4E", x"03C2", x"0AFA", x"0FD4", x"1255", x"134C", x"1397", x"13F5",
		x"1481", x"14F2", x"14B1", x"12D6", x"0EBC", x"0855", x"0076", x"F8A6",
		x"F226", x"EDCC", x"EB93", x"EACC", x"EAD2", x"EAED", x"EAFA", x"EB2F",
		x"EBCF", x"ED06", x"EF2A", x"F212", x"F576", x"F937", x"FD18", x"00E7",
		x"0439", x"0678", x"071C", x"05AF", x"01D5", x"FBF6", x"F528", x"EF3F",
		x"EC47", x"ECB0", x"EF84", x"F2B2", x"F44D", x"F36B", x"F0BE", x"EDEE",
		x"ED2C", x"EFE1", x"F5C6", x"FD49", x"047B", x"0A0B", x"0D63", x"0F18",
		x"0FCF", x"104D", x"1125", x"1271", x"13B8", x"1411", x"125E", x"0DF2",
		x"0725", x"FF47", x"F7D4", x"F1D8", x"EDFF", x"EBE4", x"EB48", x"EBA7",
		x"ECF2", x"EF11", x"F1FB", x"F511", x"F7BD", x"F915", x"F8B3", x"F6C9",
		x"F3BF", x"F0B3", x"EE16", x"EC34", x"EB36", x"EB3D", x"ED14", x"F169",
		x"F85B", x"00DF", x"08F5", x"0F36", x"1338", x"1528", x"1581", x"14BD",
		x"12CF", x"0F2C", x"0966", x"0194", x"F906", x"F182", x"ECCA", x"EAB3",
		x"EA86", x"EB28", x"EC1B", x"ECCC", x"ED6A", x"EE35", x"EF56", x"F128",
		x"F38D", x"F689", x"F9D6", x"FD37", x"0032", x"0251", x"0366", x"0352",
		x"0226", x"FFEE", x"FD01", x"F9AC", x"F677", x"F3C0", x"F1DB", x"F145",
		x"F1D4", x"F3C8", x"F6FE", x"FAF8", x"FF22", x"027E", x"0454", x"03C8",
		x"0086", x"FAD2", x"F428", x"EEEE", x"ECEB", x"EE5E", x"F20C", x"F588",
		x"F6F7", x"F57A", x"F1CD", x"EE28", x"ECDC", x"EF44", x"F46E", x"FAB2",
		x"0000", x"0317", x"03D7", x"026C", x"FF73", x"FBBF", x"F7E5", x"F447",
		x"F116", x"EEB0", x"ED07", x"EC05", x"EB65", x"EB19", x"EAE3", x"EAEB",
		x"EB68", x"EC31", x"ED7E", x"EF63", x"F19E", x"F43E", x"F6F0", x"F908",
		x"FA80", x"FB02", x"FA64", x"F8B4", x"F65A", x"F37C", x"F0B3", x"EE82",
		x"ED09", x"EC5A", x"EC75", x"ED6D", x"EF68", x"F274", x"F623", x"F9A0",
		x"FC01", x"FC48", x"F9EB", x"F59F", x"F0DF", x"ED95", x"ED4A", x"F035",
		x"F566", x"FA84", x"FD8B", x"FD1C", x"F979", x"F431", x"EF94", x"ED84",
		x"EED6", x"F326", x"F8E4", x"FED4", x"03E7", x"07AA", x"09F7", x"0B65",
		x"0C6C", x"0DA5", x"0F28", x"10DA", x"126B", x"13A8", x"148F", x"1509",
		x"1532", x"1510", x"14A3", x"13C0", x"1275", x"10A7", x"0E3F", x"0B71",
		x"085A", x"0595", x"03B0", x"02E6", x"0336", x"04F1", x"07D8", x"0B41",
		x"0E8B", x"10FF", x"12A7", x"1326", x"11B8", x"0D7C", x"0667", x"FDD0",
		x"F5BA", x"EFCF", x"EC5F", x"EAE7", x"EA82", x"EAC3", x"EC0F", x"EF24",
		x"F47F", x"FBC3", x"03C2", x"0ACA", x"0F77", x"10B6", x"0E5A", x"0907",
		x"01AD", x"F99E", x"F28C", x"EDDF", x"EC50", x"ED88", x"F039", x"F303",
		x"F51E", x"F6A9", x"F7FE", x"F992", x"FB87", x"FDFD", x"0123", x"04A5",
		x"082E", x"0B57", x"0DF1", x"0FC5", x"10E1", x"113B", x"10C3", x"0FAE",
		x"0DEE", x"0BC8", x"0971", x"070C", x"04AB", x"02C0", x"018E", x"0113",
		x"014A", x"023C", x"03FC", x"0693", x"0A14", x"0E03", x"119F", x"138E",
		x"12B6", x"0EC0", x"083B", x"0086", x"F8FA", x"F307", x"EFEC", x"EFFF",
		x"F34B", x"F967", x"0108", x"08D9", x"0F2C", x"12FB", x"142A", x"1397",
		x"12BC", x"129C", x"1370", x"148A", x"152B", x"149D", x"1330", x"114B",
		x"0F97", x"0E4E", x"0D8E", x"0CF5", x"0BD7", x"09AF", x"0615", x"011C",
		x"FB09", x"F4C3", x"EF93", x"ECCD", x"ED2B", x"F07B", x"F57B", x"FA8C",
		x"FE16", x"FF5D", x"FE6D", x"FBC3", x"F852", x"F4E2", x"F1FE", x"EFDD",
		x"EEA7", x"EEAF", x"F040", x"F356", x"F75B", x"FB89", x"FF10", x"00F1",
		x"0057", x"FCF8", x"F791", x"F1E2", x"EDFC", x"ED71", x"F02F", x"F4B8",
		x"F8B0", x"FA0A", x"F7FF", x"F37C", x"EED6", x"EC94", x"EE05", x"F2CA",
		x"F89F", x"FD8B", x"007E", x"014B", x"0052", x"FDB8", x"FA23", x"F638",
		x"F2B7", x"EFEA", x"EDE1", x"EC33", x"EAE3", x"EA11", x"E9FC", x"EA87",
		x"EB54", x"EBE0", x"EBCF", x"EB6E", x"EAE4", x"EA9A", x"EACF", x"EB6F",
		x"EC6C", x"ED7A", x"EE10", x"EE11", x"ED98", x"ECB4", x"EBD3", x"EB59",
		x"EB54", x"EB94", x"EBEF", x"EBF7", x"EBC6", x"EB92", x"EBC6", x"EC6F",
		x"ED67", x"EE1B", x"EE08", x"ED27", x"EC1F", x"EC11", x"EE53", x"F349",
		x"FA8F", x"0284", x"0967", x"0E0E", x"104D", x"1077", x"0F19", x"0C9B",
		x"095E", x"05AC", x"01CE", x"FE14", x"FAD7", x"F80D", x"F5CD", x"F3BB",
		x"F1BF", x"EFDA", x"EE0E", x"ECA9", x"EBD3", x"EB58", x"EB11", x"EAC6",
		x"EACE", x"EB1A", x"EBF4", x"ED45", x"EF11", x"F125", x"F3A6", x"F699",
		x"F986", x"FC56", x"FEAC", x"0040", x"0104", x"013C", x"0101", x"0066",
		x"FF68", x"FDBB", x"FB02", x"F762", x"F332", x"EF2F", x"ECC4", x"ECF9",
		x"F020", x"F5DF", x"FCF6", x"03FF", x"0973", x"0C5F", x"0C1E", x"08D8",
		x"0322", x"FC02", x"F4BC", x"EF4B", x"ED21", x"EF0E", x"F4A5", x"FC60",
		x"04A3", x"0BD3", x"10FE", x"13AB", x"13FF", x"129F", x"1032", x"0D50",
		x"0A76", x"0826", x"066B", x"04C3", x"02B6", x"FF96", x"FB2F", x"F5F5",
		x"F0E0", x"ED87", x"ED26", x"F01C", x"F572", x"FB89", x"007C", x"0307",
		x"02C9", x"005A", x"FCB1", x"F8D2", x"F54D", x"F31D", x"F245", x"F36E",
		x"F6A1", x"FBC1", x"0241", x"0914", x"0F12", x"12BA", x"131B", x"0F87",
		x"0882", x"FF73", x"F696", x"EFC6", x"EC34", x"EB64", x"EC41", x"ED2A",
		x"ED59", x"EC9A", x"EC10", x"ED54", x"F15E", x"F82C", x"0054", x"081B",
		x"0E0F", x"11B3", x"139C", x"1469", x"14D8", x"1510", x"152D", x"1511",
		x"14B6", x"144A", x"13A3", x"12E8", x"11D0", x"1066", x"0E3E", x"0B64",
		x"0740", x"01CA", x"FB03", x"F421", x"EEDB", x"EC7E", x"ED1C", x"EFD8",
		x"F357", x"F656", x"F83C", x"F8E8", x"F842", x"F684", x"F3FD", x"F0F8",
		x"EE07", x"EBF8", x"EC23", x"EF81", x"F5DA", x"FDFC", x"0611", x"0CCA",
		x"1192", x"13F6", x"139C", x"1038", x"0A00", x"01FC", x"F9B3", x"F27C",
		x"ED60", x"EA80", x"E9CB", x"EAFA", x"EDD4", x"F289", x"F929", x"00FC",
		x"08EE", x"0F54", x"1373", x"1519", x"1553", x"14E2", x"1412", x"12AD",
		x"1054", x"0C9A", x"079F", x"018F", x"FAEE", x"F4BA", x"EFD0", x"ECEA",
		x"EC6E", x"EE74", x"F24B", x"F768", x"FCFB", x"01F1", x"05E2", x"088C",
		x"0A23", x"0AD7", x"0B22", x"0B0C", x"0A80", x"0989", x"0837", x"0682",
		x"044D", x"017C", x"FE42", x"FA94", x"F6DA", x"F33D", x"EFFC", x"ED88",
		x"EBF9", x"EB65", x"EB5E", x"EBB1", x"EC6E", x"EDF4", x"F0FD", x"F617",
		x"FD20", x"051B", x"0C98", x"11D1", x"13A2", x"11A2", x"0C9A", x"05AC",
		x"FE59", x"F779", x"F1B6", x"ED7A", x"EB32", x"EB08", x"EC95", x"EF79",
		x"F2C3", x"F5B4", x"F76C", x"F78E", x"F620", x"F384", x"F085", x"EDC4",
		x"EC6C", x"ED4F", x"F0C3", x"F682", x"FD88", x"04AD", x"0AC1", x"0F5F",
		x"126B", x"1425", x"14D4", x"1519", x"1550", x"1508", x"13B9", x"0FD2",
		x"0946", x"00F3", x"F8A3", x"F1AD", x"ECE9", x"EA5E", x"E9D2", x"EB61",
		x"EEE9", x"F45C", x"FB8F", x"03A7", x"0B41", x"1109", x"1449", x"154C",
		x"1557", x"1517", x"14A9", x"13A8", x"118B", x"0E14", x"0977", x"03DC",
		x"FD7D", x"F6E8", x"F146", x"ED8F", x"EC44", x"ED6C", x"F0D3", x"F5A3",
		x"FAAF", x"FF19", x"01F3", x"03CD", x"0511", x"066B", x"07FF", x"09E8",
		x"0C11", x"0E54", x"10C7", x"12D1", x"146E", x"154F", x"15A4", x"15A4",
		x"1549", x"14A3", x"1397", x"1220", x"104D", x"0E8F", x"0D76", x"0D81",
		x"0EB7", x"10C6", x"12F9", x"1407", x"12DC", x"0E80", x"0778", x"FEF6",
		x"F6D0", x"F046", x"EC57", x"EB70", x"ED36", x"F128", x"F6A6", x"FD8E",
		x"053C", x"0C81", x"11BF", x"1374", x"1194", x"0CF6", x"06E5", x"00CA",
		x"FBC5", x"F874", x"F747", x"F7C5", x"F975", x"FBD5", x"FECB", x"024A",
		x"0602", x"09BD", x"0D2C", x"100B", x"1248", x"13C8", x"148A", x"14E0",
		x"153C", x"153A", x"1454", x"1187", x"0C19", x"047C", x"FC23", x"F491",
		x"EEF3", x"EBC0", x"EAC2", x"EBCA", x"EEFF", x"F466", x"FBAF", x"03FF",
		x"0BC5", x"1198", x"146E", x"1459", x"1271", x"0FA5", x"0CE1", x"0ACA",
		x"098B", x"09A1", x"0B21", x"0DDD", x"10E4", x"1321", x"1326", x"1030",
		x"0AA4", x"03BC", x"FD71", x"F906", x"F71F", x"F7C5", x"FA65", x"FE9B",
		x"0329", x"0771", x"0A6F", x"0BB2", x"0B04", x"08CB", x"054E", x"0112",
		x"FCB9", x"F955", x"F7A5", x"F858", x"FB96", x"012D", x"07FB", x"0E6C",
		x"12B5", x"139B", x"11B7", x"0E59", x"0B0C", x"092C", x"090D", x"0A71",
		x"0CE1", x"0F88", x"1209", x"13E0", x"1502", x"153B", x"14CE", x"1432",
		x"1375", x"12BD", x"11D2", x"1091", x"0EBC", x"0C47", x"0945", x"05AC",
		x"0209", x"FEA7", x"FBCC", x"F9DA", x"F8F7", x"F929", x"FA73", x"FCA3",
		x"FF9C", x"02BD", x"05C1", x"0830", x"09F1", x"0AF9", x"0B60", x"0B26",
		x"0A70", x"0934", x"072D", x"042E", x"FFB7", x"FA1C", x"F432", x"EF64",
		x"ECF6", x"ED91", x"F14C", x"F6FE", x"FCF7", x"0169", x"02D7", x"00C9",
		x"FBE7", x"F5B3", x"F02C", x"ED2F", x"ED9C", x"F107", x"F645", x"FBC0",
		x"0093", x"0426", x"06A0", x"082C", x"097B", x"0AE1", x"0C70", x"0E0C",
		x"0FA7", x"1134", x"12BD", x"13BE", x"1462", x"14C1", x"14A3", x"138E",
		x"1048", x"0A7C", x"02D4", x"FAA4", x"F376", x"EE3C", x"EB50", x"EA38",
		x"EA39", x"EAB8", x"EB56", x"EC82", x"EE0E", x"EFDF", x"F0FF", x"F0F2",
		x"EF92", x"EDF4", x"ED9D", x"F01F", x"F5A6", x"FD5E", x"050A", x"0A62",
		x"0BB4", x"0891", x"01BB", x"F97B", x"F26C", x"EE22", x"ED0F", x"EDC3",
		x"EE68", x"EE52", x"ED8C", x"ED6A", x"EF50", x"F428", x"FB5A", x"0329",
		x"09AC", x"0DB2", x"0F29", x"0E9B", x"0C74", x"091A", x"050B", x"00D7",
		x"FCD4", x"F965", x"F67C", x"F425", x"F257", x"F0C1", x"EF69", x"EE01",
		x"ECC5", x"EB9F", x"EB0F", x"EB03", x"EB83", x"EC54", x"ED51", x"EE2A",
		x"EEE5", x"EF7A", x"EF78", x"EEEE", x"EDF5", x"ECCD", x"EBC6", x"EB03",
		x"EAC0", x"EB34", x"EC4D", x"EE00", x"F025", x"F2DC", x"F5E0", x"F8B4",
		x"FA7D", x"FA82", x"F884", x"F504", x"F0E6", x"EDDB", x"ED48", x"EFDB",
		x"F4F4", x"FAE3", x"FF5E", x"0055", x"FD82", x"F7F5", x"F215", x"EE4A",
		x"EDD3", x"F09B", x"F59B", x"FB2F", x"001F", x"038F", x"05A1", x"06BF",
		x"07C4", x"0978", x"0BF6", x"0F1E", x"1206", x"138E", x"1298", x"0EA7",
		x"084A", x"00DC", x"F9E9", x"F43D", x"EFF0", x"ECDD", x"EB24", x"EA9F",
		x"EAC8", x"EB2E", x"EB92", x"EBBE", x"EBA9", x"EB62", x"EB3A", x"EB5A",
		x"EC35", x"EDA8", x"EEE0", x"EF42", x"EE5E", x"ED26", x"ECBB", x"EE72"
	);
begin
	dut: freq_demod port map(
		clk_i => clk_i,
		i_i => i_i,
		q_i => q_i,
		demod_o => demod_o
	);

	process
		variable cnt : integer range 0 to 20000 := 0;
	begin
		wait for 25 us;
		i_i <= i_vals(cnt);
		q_i <= q_vals(cnt);
		if cnt<20000 then
			cnt := cnt + 1;
		else
			cnt := 0;
		end if;
	end process;

	process
	begin
		wait for 25 us;
		clk_i <= not clk_i;
	end process;
end sim;
