-------------------------------------------------------------
-- Version declaration
--
-- Sebastien Van Cauwenberghe, ON4SEB
--
-- M17 Project
-- February 2024
-------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.math_real.all;

package version_pkg is
    constant VERSION_MAJOR: natural := 0;
    constant VERSION_MINOR: natural := 5;

end package;